* NGSPICE file created from ram_16B.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

.subckt ram_16B address[0] address[1] address[2] address[3] clk data_in[0] data_in[1]
+ data_in[2] data_in[3] data_in[4] data_in[5] data_in[6] data_in[7] data_out[0] data_out[1]
+ data_out[2] data_out[3] data_out[4] data_out[5] data_out[6] data_out[7] rd_wr vdd
+ vss
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1454__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1724__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1874__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1270_ _0799_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0985_ ram16\[0\].rb.ram1\[2\].rc.rd ram16\[0\].rb.ram1\[2\].rc.mem _0621_ _0626_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1606_ ram16\[14\].rb.ram1\[2\].rc.mem _0448_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1537_ ram16\[13\].rb.ram1\[7\].rc.mem _0403_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1468_ ram16\[11\].rb.ram1\[5\].rc.mem ram16\[11\].rb.ram1\[5\].rc.rd _0363_ _0365_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1399_ ram16\[9\].rb.ram1\[0\].rc.mem _0310_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1747__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1299__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1897__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0931__I _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0961__I0 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1203__S _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0841__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1322_ ram16\[8\].rb.ram1\[7\].rc.rd ram16\[8\].rb.ram1\[7\].rc.mem _0269_ _0271_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1253_ ram16\[6\].rb.ram1\[4\].rc.mem _0779_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1184_ _0737_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1409__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0968_ _0615_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0899_ ram16\[2\].rb.ram1\[4\].rc.rd ram16\[3\].rb.ram1\[4\].rc.rd ram16\[10\].rb.ram1\[4\].rc.rd
+ ram16\[11\].rb.ram1\[4\].rc.rd _0546_ _0522_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0943__I0 ram16\[0\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1648__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1023__S _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1912__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0836__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1871_ _0201_ clknet_leaf_51_clk ram16\[12\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1305_ _0260_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0925__I0 ram16\[2\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1236_ ram16\[5\].rb.ram1\[1\].rc.mem ram16\[5\].rb.ram1\[1\].rc.rd _0794_ _0796_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1167_ ram16\[4\].rb.ram1\[5\].rc.rd _0747_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1098_ ram16\[3\].rb.ram1\[7\].rc.rd _0696_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_22_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1808__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1021_ _0648_ ram16\[1\].rb.ram1\[2\].rc.mem _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1923_ _0253_ clknet_leaf_13_clk ram16\[14\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1854_ _0184_ clknet_leaf_15_clk ram16\[11\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1785_ _0115_ clknet_leaf_22_clk ram16\[7\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1219_ ram16\[5\].rb.ram1\[4\].rc.mem ram16\[5\].rb.ram1\[4\].rc.rd _0780_ _0785_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1242__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0426_ _0427_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1780__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1004_ _0638_ ram16\[1\].rb.ram1\[5\].rc.mem _0635_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1906_ _0236_ clknet_leaf_9_clk ram16\[14\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1837_ _0167_ clknet_leaf_3_clk ram16\[10\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1768_ _0098_ clknet_leaf_24_clk ram16\[6\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1699_ _0029_ clknet_leaf_18_clk ram16\[15\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1590__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput20 net20 data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1206__S _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0889__I2 ram16\[8\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1622_ _0406_ _0461_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1553_ ram16\[13\].rb.ram1\[3\].rc.mem _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1484_ ram16\[11\].rb.ram1\[0\].rc.mem _0793_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1390__A1 ram16\[9\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1026__S _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1133__A1 ram16\[3\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1436__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1699__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0984_ _0625_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1605_ _0620_ _0446_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1536_ ram16\[13\].rb.ram1\[7\].rc.rd _0400_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1467_ _0364_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1398_ _0728_ _0308_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1666__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1841__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1418__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0929__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1321_ _0270_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1252_ _0799_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1106__A1 ram16\[3\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1657__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1183_ _0760_ _0761_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1409__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0967_ _0613_ ram16\[0\].rb.ram1\[4\].rc.mem _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1593__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0898_ _0492_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1714__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1519_ _0393_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0943__I1 ram16\[1\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1304__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1648__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0934__I1 ram16\[1\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1639__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1214__S _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0852__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1870_ _0200_ clknet_leaf_47_clk ram16\[12\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1737__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1887__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1304_ ram16\[7\].rb.ram1\[1\].rc.mem _0790_ _0257_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0925__I1 ram16\[3\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1235_ _0795_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1166_ _0749_ _0750_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0963__S _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1097_ _0697_ _0701_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1034__S _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1557__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0907__I1 ram16\[5\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1008__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1020_ _0634_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0915__S0 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1922_ _0252_ clknet_leaf_8_clk ram16\[15\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1853_ _0183_ clknet_leaf_11_clk ram16\[11\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1784_ _0114_ clknet_leaf_23_clk ram16\[7\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0958__S _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1218_ _0784_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1149_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1902__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1539__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1242__A3 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_21_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1925__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1003_ net10 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_36_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1905_ _0235_ clknet_leaf_9_clk ram16\[14\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1836_ _0166_ clknet_leaf_32_clk ram16\[10\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1767_ _0097_ clknet_leaf_23_clk ram16\[6\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1698_ _0028_ clknet_leaf_52_clk ram16\[1\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input11_I data_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput21 net21 data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0889__I3 ram16\[9\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0860__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1621_ _0767_ _0424_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1552_ _0402_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1483_ _0357_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input3_I address[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1151__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1819_ _0149_ clknet_leaf_46_clk ram16\[9\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1390__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1217__S _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1381__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1133__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0983_ _0624_ ram16\[0\].rb.ram1\[1\].rc.mem _0621_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1604_ _0444_ _0450_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1535_ _0401_ _0404_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1466_ ram16\[11\].rb.ram1\[4\].rc.mem _0779_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1124__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1397_ _0314_ _0319_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1793__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0874__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1500__S _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0929__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1320_ _0632_ ram16\[8\].rb.ram1\[6\].rc.mem _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1251_ _0804_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1106__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1182_ ram16\[4\].rb.ram1\[1\].rc.mem _0754_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0966_ _0606_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1042__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1593__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0897_ _0512_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1518_ ram16\[12\].rb.ram1\[2\].rc.rd ram16\[12\].rb.ram1\[2\].rc.mem _0389_ _0393_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0943__I2 ram16\[8\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1449_ ram16\[10\].rb.ram1\[1\].rc.rd _0350_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1320__S _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1584__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__CLK clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0934__I2 ram16\[8\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1230__S _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1575__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1303_ _0259_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1234_ ram16\[5\].rb.ram1\[0\].rc.mem _0793_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1165_ ram16\[4\].rb.ram1\[4\].rc.mem _0741_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1096_ ram16\[3\].rb.ram1\[6\].rc.mem _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1566__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0949_ net2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1831__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1315__S _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1114__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1557__A2 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0907__I2 ram16\[12\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1225__S _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1704__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ _0251_ clknet_leaf_8_clk ram16\[15\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1852_ _0182_ clknet_leaf_25_clk ram16\[11\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1783_ _0113_ clknet_leaf_23_clk ram16\[7\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1548__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1217_ ram16\[5\].rb.ram1\[3\].rc.mem _0783_ _0780_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0974__S _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1148_ _0735_ _0698_ _0603_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1079_ _0655_ ram16\[2\].rb.ram1\[0\].rc.mem _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0948__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1242__A4 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1250__I1 ram16\[6\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1019__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1002_ _0637_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1904_ _0234_ clknet_leaf_9_clk ram16\[14\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _0165_ clknet_leaf_3_clk ram16\[10\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1766_ _0096_ clknet_leaf_19_clk ram16\[6\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0969__S _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1697_ _0027_ clknet_leaf_51_clk ram16\[1\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1503__S _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1620_ _0455_ _0460_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1223__I1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ _0617_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1482_ _0372_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1818_ _0148_ clknet_leaf_31_clk ram16\[9\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1749_ _0079_ clknet_leaf_24_clk ram16\[5\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1214__I1 ram16\[5\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1122__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_20_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1915__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_35_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0982_ net6 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1603_ ram16\[14\].rb.ram1\[4\].rc.rd _0441_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1534_ ram16\[13\].rb.ram1\[6\].rc.mem _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1465_ _0357_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1396_ ram16\[9\].rb.ram1\[2\].rc.rd _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0874__A2 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1228__S _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1250_ ram16\[6\].rb.ram1\[6\].rc.mem ram16\[6\].rb.ram1\[6\].rc.rd _0800_ _0804_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0866__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1181_ _0723_ _0752_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0965_ net9 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1042__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0896_ ram16\[0\].rb.ram1\[4\].rc.rd ram16\[1\].rb.ram1\[4\].rc.rd ram16\[8\].rb.ram1\[4\].rc.rd
+ ram16\[9\].rb.ram1\[4\].rc.rd _0514_ _0516_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0928__I0 ram16\[6\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1517_ _0392_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1448_ _0352_ _0353_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1353__I0 ram16\[8\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1379_ _0302_ _0307_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1760__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_2_2__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1344__I0 ram16\[8\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1302_ ram16\[7\].rb.ram1\[3\].rc.mem ram16\[7\].rb.ram1\[3\].rc.rd _0257_ _0259_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0925__I3 ram16\[11\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1233_ _0772_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1335__I0 ram16\[8\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1164_ _0709_ _0738_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1095_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0948_ net11 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0879_ _0520_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1326__I0 ram16\[8\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1331__S _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1920_ _0250_ clknet_leaf_8_clk ram16\[15\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1851_ _0181_ clknet_leaf_15_clk ram16\[11\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1782_ _0112_ clknet_leaf_19_clk ram16\[7\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1181__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1216_ net8 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1147_ _0494_ _0491_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1078_ _0671_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1326__S _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1061__S _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1236__S _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1001_ ram16\[1\].rb.ram1\[7\].rc.rd ram16\[1\].rb.ram1\[7\].rc.mem _0635_ _0637_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1821__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1903_ _0233_ clknet_leaf_9_clk ram16\[14\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1834_ _0164_ clknet_leaf_31_clk ram16\[10\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1765_ _0095_ clknet_leaf_23_clk ram16\[6\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1696_ _0026_ clknet_leaf_48_clk ram16\[1\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0985__S _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1056__S _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1448__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1844__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_9_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1550_ _0399_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ ram16\[11\].rb.ram1\[2\].rc.mem ram16\[11\].rb.ram1\[2\].rc.rd _0368_ _0372_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1136__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1611__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1817_ _0147_ clknet_leaf_34_clk ram16\[9\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1717__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1748_ _0078_ clknet_leaf_6_clk ram16\[4\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1679_ _0009_ clknet_leaf_4_clk ram16\[0\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1867__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1514__S _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0981_ _0623_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _0447_ _0449_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1533_ _0402_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1464_ _0362_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1395_ _0291_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_30_clk clknet_2_1__leaf_clk clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1587__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1509__S _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1308__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1244__S _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1180_ _0755_ _0759_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0945__S0 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0964_ _0612_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0895_ _0503_ _0551_ _0510_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1516_ _0652_ ram16\[12\].rb.ram1\[1\].rc.mem _0389_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1447_ ram16\[10\].rb.ram1\[0\].rc.mem _0342_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1378_ ram16\[9\].rb.ram1\[5\].rc.rd _0303_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0936__S0 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0993__S _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1905__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1329__S _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0919__I1 ram16\[7\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1128__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1032__I0 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1301_ _0258_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1232_ net5 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1163_ _0742_ _0748_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1094_ _0515_ _0698_ _0604_ _0694_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_92_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0947_ _0593_ _0595_ _0597_ _0599_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0878_ _0492_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1023__I0 ram16\[1\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1326__I1 ram16\[8\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1411__I _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1190__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1850_ _0180_ clknet_leaf_26_clk ram16\[11\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1781_ _0111_ clknet_leaf_24_clk ram16\[7\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1750__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1181__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1215_ _0782_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1146_ _0505_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1077_ _0686_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1172__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1342__S _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1141__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1773__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1000_ _0636_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1051__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1902_ _0232_ clknet_leaf_13_clk ram16\[14\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1833_ _0163_ clknet_leaf_32_clk ram16\[10\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1764_ _0094_ clknet_leaf_7_clk ram16\[5\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1695_ _0025_ clknet_2_0__leaf_clk ram16\[1\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1129_ _0723_ _0714_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1796__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1090__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1393__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1072__S _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ _0371_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1136__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1816_ _0146_ clknet_leaf_31_clk ram16\[9\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1747_ _0077_ clknet_leaf_43_clk ram16\[3\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1375__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1678_ _0008_ clknet_leaf_6_clk ram16\[0\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0886__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1067__S _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1366__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1811__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1118__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0980_ ram16\[0\].rb.ram1\[3\].rc.rd ram16\[0\].rb.ram1\[3\].rc.mem _0621_ _0623_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1601_ ram16\[14\].rb.ram1\[3\].rc.mem _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1532_ _0495_ _0294_ _0525_ _0295_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1463_ ram16\[11\].rb.ram1\[6\].rc.mem ram16\[11\].rb.ram1\[6\].rc.rd _0358_ _0362_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1109__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I address[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ _0316_ _0317_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1596__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_8_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1587__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1525__S _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1707__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0873__I1 ram16\[1\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1857__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0963_ ram16\[0\].rb.ram1\[6\].rc.rd ram16\[0\].rb.ram1\[6\].rc.mem _0607_ _0612_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_0894_ ram16\[4\].rb.ram1\[4\].rc.rd ram16\[5\].rb.ram1\[4\].rc.rd ram16\[12\].rb.ram1\[4\].rc.rd
+ ram16\[13\].rb.ram1\[4\].rc.rd _0540_ _0506_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1515_ _0391_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1446_ _0728_ _0340_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1377_ _0305_ _0306_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1569__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1319__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0863__S0 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1255__S _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1300_ ram16\[7\].rb.ram1\[2\].rc.mem _0786_ _0257_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1231_ _0792_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1162_ ram16\[4\].rb.ram1\[6\].rc.rd _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1093_ net3 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0946_ _0555_ _0598_ _0572_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1271__I1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0877_ _0529_ _0531_ _0533_ _0535_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1429_ _0713_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1262__I1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1780_ _0110_ clknet_leaf_12_clk ram16\[6\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1253__I1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1049__I _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0888__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_33_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1214_ ram16\[5\].rb.ram1\[5\].rc.mem ram16\[5\].rb.ram1\[5\].rc.rd _0780_ _0782_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_48_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1145_ _0730_ _0734_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1076_ ram16\[2\].rb.ram1\[2\].rc.rd ram16\[2\].rb.ram1\[2\].rc.mem _0682_ _0686_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0999__S _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1244__I1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0929_ _0519_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1918__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1901_ _0231_ clknet_leaf_9_clk ram16\[14\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1832_ _0162_ clknet_leaf_32_clk ram16\[10\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1763_ _0093_ clknet_leaf_30_clk ram16\[4\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1694_ _0024_ clknet_leaf_45_clk ram16\[1\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0985__I0 ram16\[0\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1128_ net6 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1059_ _0676_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1090__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1217__I1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput14 net14 data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1353__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1152__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1605__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1208__I1 ram16\[5\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1890__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0967__I0 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1815_ _0145_ clknet_leaf_34_clk ram16\[9\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1746_ _0076_ clknet_leaf_0_clk ram16\[4\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1677_ _0007_ clknet_leaf_29_clk ram16\[0\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0886__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1763__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1083__S _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1600_ _0434_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1357__A3 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1531_ _0600_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1462_ _0361_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1786__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1393_ ram16\[9\].rb.ram1\[1\].rc.mem _0310_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1520__I _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1045__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1729_ _0059_ clknet_leaf_2_clk ram16\[3\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1430__I _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1347__I0 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0873__I2 ram16\[8\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0962_ _0611_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0893_ _0536_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1514_ ram16\[12\].rb.ram1\[3\].rc.rd ram16\[12\].rb.ram1\[3\].rc.mem _0389_ _0391_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1338__I0 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1445_ _0346_ _0351_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1376_ ram16\[9\].rb.ram1\[4\].rc.mem _0297_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1451__S _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1329__I0 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0863__S1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1193__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0940__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1230_ ram16\[5\].rb.ram1\[2\].rc.mem ram16\[5\].rb.ram1\[2\].rc.rd _0787_ _0792_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1161_ _0737_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1271__S _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1092_ _0692_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1824__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0945_ ram16\[2\].rb.ram1\[0\].rc.rd ram16\[3\].rb.ram1\[0\].rc.rd ram16\[10\].rb.ram1\[0\].rc.rd
+ ram16\[11\].rb.ram1\[0\].rc.rd _0504_ _0570_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0876_ _0519_ _0534_ _0526_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1428_ _0325_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1359_ _0692_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0922__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1847__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1266__S _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0913__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1213_ _0781_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1144_ ram16\[3\].rb.ram1\[0\].rc.rd _0726_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1075_ _0685_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0928_ ram16\[6\].rb.ram1\[1\].rc.rd ram16\[7\].rb.ram1\[1\].rc.rd ram16\[14\].rb.ram1\[1\].rc.rd
+ ram16\[15\].rb.ram1\[1\].rc.rd _0521_ _0558_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0859_ _0492_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0904__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1632__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1613__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1900_ _0230_ clknet_leaf_19_clk ram16\[14\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1623__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1831_ _0161_ clknet_leaf_32_clk ram16\[10\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1762_ _0092_ clknet_leaf_7_clk ram16\[5\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1387__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ _0023_ clknet_leaf_48_clk ram16\[1\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1139__A1 ram16\[3\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1127_ _0717_ _0722_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1058_ ram16\[2\].rb.ram1\[6\].rc.rd ram16\[2\].rb.ram1\[6\].rc.mem _0672_ _0676_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1614__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1378__A1 ram16\[9\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1692__CLK clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput15 net15 data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1605__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_51_clk clknet_2_0__leaf_clk clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_32_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1369__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_47_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_42_clk clknet_2_1__leaf_clk clknet_leaf_42_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1814_ _0144_ clknet_leaf_43_clk ram16\[9\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1745_ _0075_ clknet_leaf_0_clk ram16\[4\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1676_ _0006_ clknet_leaf_4_clk ram16\[0\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1532__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1908__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1599__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_clk clknet_2_1__leaf_clk clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1428__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0885__I0 ram16\[2\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk clknet_leaf_24_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1461_ ram16\[11\].rb.ram1\[5\].rc.mem _0776_ _0358_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1392_ _0723_ _0308_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_clk clknet_2_2__leaf_clk clknet_leaf_15_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1728_ _0058_ clknet_leaf_2_clk ram16\[3\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1659_ _0627_ _0473_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0939__S0 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0961_ _0610_ ram16\[0\].rb.ram1\[5\].rc.mem _0607_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0892_ ram16\[6\].rb.ram1\[4\].rc.rd ram16\[7\].rb.ram1\[4\].rc.rd ram16\[14\].rb.ram1\[4\].rc.rd
+ ram16\[15\].rb.ram1\[4\].rc.rd _0537_ _0498_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__1753__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ _0390_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_4_clk clknet_2_2__leaf_clk clknet_leaf_4_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1444_ ram16\[10\].rb.ram1\[2\].rc.rd _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1375_ _0709_ _0292_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1026__I0 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1017__I0 ram16\[1\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1193__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0940__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1160_ _0745_ _0746_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1091_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0944_ _0545_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0875_ ram16\[2\].rb.ram1\[6\].rc.rd ram16\[3\].rb.ram1\[6\].rc.rd ram16\[10\].rb.ram1\[6\].rc.rd
+ ram16\[11\].rb.ram1\[6\].rc.rd _0521_ _0522_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1427_ _0334_ _0339_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1358_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1261__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1289_ _0826_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1171__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1346__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0913__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1282__S _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1212_ ram16\[5\].rb.ram1\[4\].rc.mem _0779_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1143_ _0733_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1074_ _0652_ ram16\[2\].rb.ram1\[1\].rc.mem _0682_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0927_ _0575_ _0577_ _0579_ _0581_ net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1457__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0858_ _0512_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0904__A2 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0840__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1396__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1814__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1148__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1830_ _0160_ clknet_leaf_43_clk ram16\[10\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1761_ _0091_ clknet_leaf_7_clk ram16\[5\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1387__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1692_ _0022_ clknet_leaf_39_clk ram16\[1\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1139__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1126_ ram16\[3\].rb.ram1\[3\].rc.rd _0707_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1057_ _0675_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1090__A4 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1378__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1837__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput16 net16 data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1369__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1813_ _0143_ clknet_leaf_34_clk ram16\[9\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1744_ _0074_ clknet_leaf_1_clk ram16\[4\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1675_ _0005_ clknet_leaf_30_clk ram16\[0\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1470__S _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0894__I1 ram16\[5\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1109_ _0709_ _0696_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1599__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1460_ _0360_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1391_ _0311_ _0315_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1682__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1727_ _0057_ clknet_leaf_2_clk ram16\[3\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1658_ _0479_ _0484_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1589_ _0439_ _0440_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0939__S1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_31_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_46_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0875__S0 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0960_ net10 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0891_ _0539_ _0542_ _0544_ _0548_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1512_ _0648_ ram16\[12\].rb.ram1\[2\].rc.mem _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1443_ _0325_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1374_ _0298_ _0304_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0872__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0857__S0 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1090_ _0515_ _0693_ _0604_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_80_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1720__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0839__S0 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0943_ ram16\[0\].rb.ram1\[0\].rc.rd ram16\[1\].rb.ram1\[0\].rc.rd ram16\[8\].rb.ram1\[0\].rc.rd
+ ram16\[9\].rb.ram1\[0\].rc.rd _0566_ _0567_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0874_ _0512_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1870__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1426_ ram16\[10\].rb.ram1\[5\].rc.rd _0335_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1357_ _0289_ _0290_ _0693_ _0662_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1288_ ram16\[7\].rb.ram1\[6\].rc.mem ram16\[7\].rb.ram1\[6\].rc.rd _0822_ _0826_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1486__I1 ram16\[11\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1893__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1211_ _0772_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1142_ _0732_ ram16\[2\].rb.ram1\[7\].rc.mem _0687_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1073_ _0684_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__I1 ram16\[11\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0926_ _0555_ _0580_ _0572_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0857_ ram16\[0\].rb.ram1\[7\].rc.rd ram16\[1\].rb.ram1\[7\].rc.rd ram16\[8\].rb.ram1\[7\].rc.rd
+ ram16\[9\].rb.ram1\[7\].rc.rd _0514_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1409_ _0692_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1766__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0912__I0 ram16\[2\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1468__I1 ram16\[11\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0840__A2 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0903__I0 ram16\[6\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1459__I1 ram16\[11\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1760_ _0090_ clknet_leaf_5_clk ram16\[5\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1691_ _0021_ clknet_leaf_46_clk ram16\[1\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1293__S _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1789__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1125_ _0720_ _0721_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1056_ _0638_ ram16\[2\].rb.ram1\[5\].rc.mem _0672_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1468__S _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1889_ _0219_ clknet_leaf_6_clk ram16\[13\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0909_ _0561_ _0563_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput17 net17 data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1288__S _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1812_ _0142_ clknet_leaf_51_clk ram16\[8\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1087__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1743_ _0073_ clknet_leaf_0_clk ram16\[4\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1674_ _0004_ clknet_leaf_17_clk ram16\[0\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1532__A3 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0894__I2 ram16\[12\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1108_ net9 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1039_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_5_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1390_ ram16\[9\].rb.ram1\[3\].rc.rd _0303_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1827__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1726_ _0056_ clknet_leaf_44_clk ram16\[3\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1657_ ram16\[15\].rb.ram1\[2\].rc.rd _0480_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1588_ ram16\[14\].rb.ram1\[5\].rc.mem _0435_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1481__S _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1441__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0875__S1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_0__f_clk clknet_0_clk clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0890_ _0545_ _0547_ _0526_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1511_ _0378_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1442_ _0348_ _0349_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1373_ ram16\[9\].rb.ram1\[6\].rc.rd _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1120__A1 ram16\[3\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1423__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0857__S1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1187__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1275__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1709_ _0039_ clknet_leaf_50_clk ram16\[2\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1662__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1414__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1672__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1102__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0839__S1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0942_ _0561_ _0594_ _0564_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1405__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0873_ ram16\[0\].rb.ram1\[6\].rc.rd ram16\[1\].rb.ram1\[6\].rc.rd ram16\[8\].rb.ram1\[6\].rc.rd
+ ram16\[9\].rb.ram1\[6\].rc.rd _0514_ _0516_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_45_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1425_ _0337_ _0338_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1356_ _0601_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1287_ _0825_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__CLK clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0902__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1643__I _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1210_ net9 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1141_ net12 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1072_ ram16\[2\].rb.ram1\[3\].rc.rd ram16\[2\].rb.ram1\[3\].rc.mem _0682_ _0684_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1626__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0925_ ram16\[2\].rb.ram1\[2\].rc.rd ram16\[3\].rb.ram1\[2\].rc.rd ram16\[10\].rb.ram1\[2\].rc.rd
+ ram16\[11\].rb.ram1\[2\].rc.rd _0546_ _0570_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0856_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1562__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1408_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1339_ _0280_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1617__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1710__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1608__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1860__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1690_ _0020_ clknet_leaf_39_clk ram16\[1\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1124_ ram16\[3\].rb.ram1\[2\].rc.mem _0716_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1055_ _0674_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_45_clk clknet_2_0__leaf_clk clknet_leaf_45_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1083__I0 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1888_ _0218_ clknet_leaf_7_clk ram16\[13\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0908_ _0509_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0839_ ram16\[6\].rb.ram1\[7\].rc.rd ram16\[7\].rb.ram1\[7\].rc.rd ram16\[14\].rb.ram1\[7\].rc.rd
+ ram16\[15\].rb.ram1\[7\].rc.rd _0495_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__1484__S _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1733__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1883__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_36_clk clknet_2_1__leaf_clk clknet_leaf_36_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1074__I0 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_27_clk clknet_2_3__leaf_clk clknet_leaf_27_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1811_ _0141_ clknet_leaf_19_clk ram16\[7\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1065__I0 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1756__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1742_ _0072_ clknet_leaf_4_clk ram16\[4\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1673_ _0003_ clknet_leaf_39_clk ram16\[0\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1532__A4 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_clk clknet_2_3__leaf_clk clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1107_ _0701_ _0708_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1038_ _0496_ net13 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1479__S _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0910__I _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0885__I3 ram16\[11\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1779__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1047__I0 ram16\[1\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1651__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ _0055_ clknet_leaf_45_clk ram16\[3\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1656_ _0482_ _0483_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1587_ _0610_ _0432_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1921__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0905__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1510_ _0388_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1441_ ram16\[10\].rb.ram1\[1\].rc.mem _0342_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1372_ _0291_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_4_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1120__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1187__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1708_ _0038_ clknet_leaf_39_clk ram16\[2\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1639_ ram16\[15\].rb.ram1\[5\].rc.rd _0465_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0870__A1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1817__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1102__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0941_ ram16\[4\].rb.ram1\[0\].rc.rd ram16\[5\].rb.ram1\[0\].rc.rd ram16\[12\].rb.ram1\[0\].rc.rd
+ ram16\[13\].rb.ram1\[0\].rc.rd _0585_ _0562_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0872_ _0503_ _0530_ _0510_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1424_ ram16\[10\].rb.ram1\[4\].rc.mem _0329_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1355_ _0670_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_68_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1286_ ram16\[7\].rb.ram1\[5\].rc.mem _0776_ _0822_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1399__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1571__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1140_ _0725_ _0731_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0921__I2 ram16\[12\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1071_ _0683_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0924_ _0512_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0855_ _0496_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1562__A2 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1407_ _0585_ _0294_ _0693_ _0662_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_84_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1338_ _0648_ ram16\[8\].rb.ram1\[2\].rc.mem _0279_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1269_ _0814_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1010__S _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1553__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_44_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1685__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1123_ _0719_ _0714_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1054_ ram16\[2\].rb.ram1\[7\].rc.rd ram16\[2\].rb.ram1\[7\].rc.mem _0672_ _0674_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0907_ ram16\[4\].rb.ram1\[3\].rc.rd ram16\[5\].rb.ram1\[3\].rc.rd ram16\[12\].rb.ram1\[3\].rc.rd
+ ram16\[13\].rb.ram1\[3\].rc.rd _0540_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1887_ _0217_ clknet_leaf_6_clk ram16\[13\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0838_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput19 net19 data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0908__I _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1474__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0896__S0 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1810_ _0140_ clknet_leaf_52_clk ram16\[8\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1741_ _0071_ clknet_leaf_0_clk ram16\[4\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1672_ _0002_ clknet_leaf_30_clk ram16\[0\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1106_ ram16\[3\].rb.ram1\[6\].rc.rd _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1037_ _0584_ _0601_ _0524_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1700__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1850__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1295__I1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1286__I1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0869__S0 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1723__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1435__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1873__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ _0054_ clknet_leaf_33_clk ram16\[3\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1655_ ram16\[15\].rb.ram1\[1\].rc.mem _0475_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1586_ _0437_ _0438_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1201__I1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1746__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1417__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1896__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0831__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1440_ _0723_ _0340_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1371_ _0301_ _0302_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1707_ _0037_ clknet_leaf_47_clk ram16\[2\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1638_ _0470_ _0471_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1569_ ram16\[13\].rb.ram1\[0\].rc.mem _0416_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0916__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0870__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0940_ _0519_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0871_ ram16\[4\].rb.ram1\[6\].rc.rd ram16\[5\].rb.ram1\[6\].rc.rd ram16\[12\].rb.ram1\[6\].rc.rd
+ ram16\[13\].rb.ram1\[6\].rc.rd _0504_ _0506_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1911__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1423_ _0709_ _0326_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1354_ _0288_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1285_ _0824_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1580__A3 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1340__I0 ram16\[8\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1096__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_3_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1070_ _0648_ ram16\[2\].rb.ram1\[2\].rc.mem _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1331__I0 ram16\[8\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0923_ ram16\[0\].rb.ram1\[2\].rc.rd ram16\[1\].rb.ram1\[2\].rc.rd ram16\[8\].rb.ram1\[2\].rc.rd
+ ram16\[9\].rb.ram1\[2\].rc.rd _0566_ _0567_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0854_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1406_ _0321_ _0324_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1337_ _0268_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1268_ ram16\[6\].rb.ram1\[2\].rc.mem ram16\[6\].rb.ram1\[2\].rc.rd _0810_ _0814_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0912__I3 ram16\[11\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1199_ _0670_ _0491_ _0508_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__1322__I0 ram16\[8\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1807__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1498__S _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1201__S _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1122_ net7 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1053_ _0673_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0906_ _0505_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1886_ _0216_ clknet_leaf_4_clk ram16\[13\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0837_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1021__S _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0834__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0896__S1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1740_ _0070_ clknet_leaf_27_clk ram16\[4\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1671_ _0001_ clknet_leaf_42_clk ram16\[0\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I data_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1105_ _0695_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1150__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1036_ net12 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1453__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1869_ _0199_ clknet_leaf_50_clk ram16\[12\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_43_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1516__I0 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1444__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1675__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1507__I0 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1435__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0869__S1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1199__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1723_ _0053_ clknet_leaf_44_clk ram16\[3\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1395__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0946__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1654_ _0624_ _0473_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1585_ ram16\[14\].rb.ram1\[7\].rc.mem _0435_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1123__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1019_ net7 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1426__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1698__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0937__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1362__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1417__A2 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1370_ ram16\[9\].rb.ram1\[5\].rc.mem _0297_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1840__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1706_ _0036_ clknet_leaf_36_clk ram16\[2\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1637_ ram16\[15\].rb.ram1\[4\].rc.mem _0667_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1568_ _0627_ _0414_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ _0382_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1713__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0941__S0 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1003__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0842__I _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0870_ _0493_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1422_ _0330_ _0336_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1353_ ram16\[8\].rb.ram1\[0\].rc.rd ram16\[8\].rb.ram1\[0\].rc.mem _0284_ _0288_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1284_ ram16\[7\].rb.ram1\[7\].rc.mem ram16\[7\].rb.ram1\[7\].rc.rd _0822_ _0824_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1629__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0932__S0 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0999_ _0632_ ram16\[1\].rb.ram1\[6\].rc.mem _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1580__A4 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0915__I1 ram16\[1\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0923__S0 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1493__I _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1331__I1 ram16\[8\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1759__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0922_ _0561_ _0576_ _0564_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0853_ net1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1405_ ram16\[9\].rb.ram1\[0\].rc.rd _0318_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1336_ _0278_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 address[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1267_ _0813_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_48_clk clknet_2_0__leaf_clk clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1198_ _0735_ _0603_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1578__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1010__I0 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_39_clk clknet_2_1__leaf_clk clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1313__I1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1901__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_0_clk_I clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1121_ _0711_ _0718_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1052_ _0632_ ram16\[2\].rb.ram1\[6\].rc.mem _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1304__I1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0905_ _0502_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1885_ _0215_ clknet_leaf_7_clk ram16\[13\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0836_ net4 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1319_ _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1924__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_2_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1302__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1101__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1212__S _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0850__I _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1670_ _0000_ clknet_leaf_42_clk ram16\[0\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1525__I1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1104_ _0705_ _0706_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1150__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1035_ _0658_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0961__S _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ _0198_ clknet_2_1__leaf_clk ram16\[12\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1799_ _0129_ clknet_leaf_38_clk ram16\[8\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1032__S _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0845__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1722_ _0052_ clknet_leaf_33_clk ram16\[3\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1653_ _0476_ _0481_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1584_ ram16\[14\].rb.ram1\[7\].rc.rd _0432_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0956__S _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1123__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1018_ _0647_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1792__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1050__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_42_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1705_ _0035_ clknet_leaf_40_clk ram16\[2\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1636_ _0613_ _0664_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1567_ _0420_ _0425_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ _0638_ ram16\[12\].rb.ram1\[5\].rc.mem _0379_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1280__A1 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0941__S1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1421_ ram16\[10\].rb.ram1\[6\].rc.rd _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1352_ _0287_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1283_ _0823_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1688__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0932__S1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0998_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1619_ ram16\[14\].rb.ram1\[1\].rc.rd _0456_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1317__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0915__I2 ram16\[8\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0923__S1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1830__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1014__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1492__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0853__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0921_ ram16\[4\].rb.ram1\[2\].rc.rd ram16\[5\].rb.ram1\[2\].rc.rd ram16\[12\].rb.ram1\[2\].rc.rd
+ ram16\[13\].rb.ram1\[2\].rc.rd _0540_ _0562_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0852_ _0502_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1404_ _0323_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1335_ ram16\[8\].rb.ram1\[4\].rc.rd ram16\[8\].rb.ram1\[4\].rc.mem _0274_ _0278_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput2 address[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1266_ ram16\[6\].rb.ram1\[1\].rc.mem _0790_ _0810_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1197_ net11 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1853__CLK clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1009__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0848__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1120_ ram16\[3\].rb.ram1\[4\].rc.rd _0707_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1051_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1726__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0899__S0 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1876__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1884_ _0214_ clknet_leaf_28_clk ram16\[13\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0904_ _0536_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0835_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1240__I1 ram16\[5\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1318_ _0602_ _0267_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1249_ _0803_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1899__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1470__I1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1103_ ram16\[3\].rb.ram1\[5\].rc.mem _0700_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1403__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1034_ ram16\[1\].rb.ram1\[1\].rc.rd ram16\[1\].rb.ram1\[1\].rc.mem _0656_ _0658_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1610__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1461__I1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _0197_ clknet_leaf_47_clk ram16\[12\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1798_ _0128_ clknet_leaf_41_clk ram16\[8\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0972__I0 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1313__S _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0951__I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1668__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1223__S _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0861__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1199__A3 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1721_ _0051_ clknet_leaf_33_clk ram16\[3\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1652_ ram16\[15\].rb.ram1\[3\].rc.rd _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_2_1__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__CLK clknet_leaf_21_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_1_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1583_ _0433_ _0436_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1659__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0972__S _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1017_ ram16\[1\].rb.ram1\[4\].rc.rd ram16\[1\].rb.ram1\[4\].rc.mem _0642_ _0647_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1919_ _0249_ clknet_leaf_8_clk ram16\[15\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0945__I0 ram16\[2\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1362__A3 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0936__I0 ram16\[2\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0856__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0034_ clknet_leaf_35_clk ram16\[2\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1635_ _0464_ _0469_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1566_ ram16\[13\].rb.ram1\[2\].rc.rd _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0967__S _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1497_ _0381_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1280__A2 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1099__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ _0325_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1351_ ram16\[7\].rb.ram1\[7\].rc.mem _0818_ _0262_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1282_ ram16\[7\].rb.ram1\[6\].rc.mem _0770_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1210__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0997_ _0513_ _0501_ _0633_ _0605_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_118_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1618_ _0458_ _0459_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1549_ _0408_ _0413_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1573__I0 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0915__I3 ram16\[9\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1782__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_41_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0920_ _0536_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1030__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0851_ _0503_ _0507_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1403_ _0732_ ram16\[8\].rb.ram1\[7\].rc.mem _0284_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1334_ _0277_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1265_ _0812_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1205__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 address[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1196_ _0765_ _0769_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0980__S _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1115__I _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1678__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1529__A3 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1025__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1050_ _0670_ _0491_ _0633_ _0605_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__0864__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0899__S1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0903_ ram16\[6\].rb.ram1\[3\].rc.rd ram16\[7\].rb.ram1\[3\].rc.rd ram16\[14\].rb.ram1\[3\].rc.rd
+ ram16\[15\].rb.ram1\[3\].rc.rd _0537_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1883_ _0213_ clknet_leaf_14_clk ram16\[13\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0834_ net1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0900__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1317_ _0496_ net13 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1248_ ram16\[6\].rb.ram1\[5\].rc.mem _0776_ _0800_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1179_ ram16\[4\].rb.ram1\[3\].rc.rd _0747_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1820__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1392__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0949__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1144__A1 ram16\[3\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1447__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1102_ _0704_ _0696_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1033_ _0657_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1843__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1438__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1610__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1866_ _0196_ clknet_leaf_36_clk ram16\[12\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1797_ _0127_ clknet_leaf_34_clk ram16\[8\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1429__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1601__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1716__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1668__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1199__A4 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1720_ _0050_ clknet_leaf_33_clk ram16\[3\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1651_ _0663_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1582_ ram16\[14\].rb.ram1\[6\].rc.mem _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1659__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I data_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1016_ _0646_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1918_ _0248_ clknet_leaf_14_clk ram16\[15\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1739__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1849_ _0179_ clknet_leaf_25_clk ram16\[11\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1889__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0945__I1 ram16\[3\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1362__A4 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1324__S _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1050__A3 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0936__I1 ram16\[3\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1234__S _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk clknet_leaf_11_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__1577__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1703_ _0033_ clknet_leaf_36_clk ram16\[2\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1634_ ram16\[15\].rb.ram1\[6\].rc.rd _0465_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1565_ _0399_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1496_ ram16\[12\].rb.ram1\[7\].rc.rd ram16\[12\].rb.ram1\[7\].rc.mem _0379_ _0381_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0983__S _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0863__I0 ram16\[2\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1568__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1054__S _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1904__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_0_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1350_ _0286_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1281_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0996_ _0508_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1617_ ram16\[14\].rb.ram1\[0\].rc.mem _0448_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0978__S _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1548_ ram16\[13\].rb.ram1\[5\].rc.rd _0409_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1479_ ram16\[11\].rb.ram1\[1\].rc.mem _0790_ _0368_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1512__S _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0850_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1402_ _0317_ _0322_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1333_ _0645_ ram16\[8\].rb.ram1\[3\].rc.mem _0274_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1264_ ram16\[6\].rb.ram1\[3\].rc.mem ram16\[6\].rb.ram1\[3\].rc.rd _0810_ _0812_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput4 address[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_1195_ ram16\[4\].rb.ram1\[0\].rc.rd _0762_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1__f_clk clknet_0_clk clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1221__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0979_ _0622_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1507__S _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1162__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1041__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0902_ _0497_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1882_ _0212_ clknet_leaf_28_clk ram16\[13\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0833_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1316_ _0266_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1216__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1153__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1247_ _0802_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1178_ _0757_ _0758_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0991__S _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_40_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1392__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1144__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0965__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1383__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1036__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1101_ net10 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1032_ _0655_ ram16\[1\].rb.ram1\[0\].rc.mem _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1865_ _0195_ clknet_leaf_40_clk ram16\[12\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1796_ _0126_ clknet_leaf_10_clk ram16\[7\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1126__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0909__B _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0876__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ _0478_ _0479_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1581_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1810__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0867__A1 _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1015_ _0645_ ram16\[1\].rb.ram1\[3\].rc.mem _0642_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ _0247_ clknet_leaf_8_clk ram16\[15\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1848_ _0178_ clknet_leaf_26_clk ram16\[11\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1779_ _0109_ clknet_leaf_17_clk ram16\[5\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0858__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1340__S _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1833__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1250__S _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1702_ _0032_ clknet_leaf_41_clk ram16\[2\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1633_ _0467_ _0468_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0880__S0 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1564_ _0422_ _0423_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1495_ _0380_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0863__I1 ram16\[3\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1856__CLK clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1568__A2 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0871__S0 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1335__S _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1070__S _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0922__B _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1280_ _0771_ _0660_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1044__I _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0995_ net11 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1616_ _0627_ _0446_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _0411_ _0412_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1478_ _0370_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1238__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1065__S _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1039__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1401_ ram16\[9\].rb.ram1\[1\].rc.rd _0318_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1332_ _0276_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1263_ _0811_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput5 data_in[0] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1194_ _0703_ _0768_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1502__I _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0978_ _0620_ ram16\[0\].rb.ram1\[2\].rc.mem _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0989__S _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1631__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1234__I1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0993__I0 ram16\[0\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1523__S _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1881_ _0211_ clknet_leaf_29_clk ram16\[13\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0901_ _0550_ _0552_ _0554_ _0557_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0832_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1225__I1 ram16\[5\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1315_ ram16\[7\].rb.ram1\[0\].rc.mem ram16\[7\].rb.ram1\[0\].rc.rd _0262_ _0266_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1246_ ram16\[6\].rb.ram1\[7\].rc.mem ram16\[6\].rb.ram1\[7\].rc.rd _0800_ _0802_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1232__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1177_ ram16\[4\].rb.ram1\[2\].rc.mem _0754_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1518__S _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1253__S _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1100_ _0702_ _0703_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1031_ _0634_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1864_ _0194_ clknet_leaf_36_clk ram16\[12\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1795_ _0125_ clknet_leaf_19_clk ram16\[6\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1227__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1229_ _0791_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1338__S _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0976__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1762__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1600__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1248__S _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1580_ _0289_ _0290_ _0693_ _0295_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_4_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1014_ net8 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1916_ _0246_ clknet_leaf_18_clk ram16\[15\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1847_ _0177_ clknet_leaf_26_clk ram16\[11\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1778_ _0108_ clknet_leaf_12_clk ram16\[6\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0858__A2 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1420__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0936__I3 ram16\[11\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1577__A3 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1701_ _0031_ clknet_leaf_35_clk ram16\[2\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1632_ ram16\[15\].rb.ram1\[5\].rc.mem _0667_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0880__S1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1563_ ram16\[13\].rb.ram1\[1\].rc.mem _0416_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1494_ _0632_ ram16\[12\].rb.ram1\[6\].rc.mem _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0871__S1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1351__S _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1500__I0 ram16\[12\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1800__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1060__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0994_ _0631_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1615_ _0452_ _0457_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1546_ ram16\[13\].rb.ram1\[4\].rc.mem _0403_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1477_ ram16\[11\].rb.ram1\[3\].rc.mem ram16\[11\].rb.ram1\[3\].rc.rd _0368_ _0370_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1823__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1238__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0997__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1081__S _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0933__B _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1401__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1400_ _0320_ _0321_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1331_ ram16\[8\].rb.ram1\[5\].rc.rd ram16\[8\].rb.ram1\[5\].rc.mem _0274_ _0276_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1262_ ram16\[6\].rb.ram1\[2\].rc.mem _0786_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1846__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 data_in[1] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1193_ _0767_ _0726_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0977_ _0606_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1529_ _0289_ _0290_ _0633_ _0662_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1719__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1076__S _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1869__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0900_ _0555_ _0556_ _0526_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _0210_ clknet_leaf_28_clk ram16\[13\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0831_ net2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1386__A1 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1314_ _0265_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1245_ _0801_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1176_ _0719_ _0752_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1129__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_50_clk clknet_2_0__leaf_clk clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1691__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1030_ net5 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_clk clknet_2_1__leaf_clk clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1863_ _0193_ clknet_leaf_36_clk ram16\[12\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1794_ _0124_ clknet_leaf_10_clk ram16\[7\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1359__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1531__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1243__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1228_ ram16\[5\].rb.ram1\[1\].rc.mem _0790_ _0787_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1159_ ram16\[4\].rb.ram1\[5\].rc.mem _0741_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_32_clk clknet_2_1__leaf_clk clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1070__I0 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk clknet_leaf_23_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1328__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1061__I0 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1264__S _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1013_ _0644_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0875__I0 ram16\[2\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1915_ _0245_ clknet_leaf_14_clk ram16\[15\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_14_clk clknet_2_2__leaf_clk clknet_leaf_14_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__0851__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _0176_ clknet_leaf_17_clk ram16\[11\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1777_ _0107_ clknet_leaf_12_clk ram16\[6\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1052__I0 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I data_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1349__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0987__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1259__S _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1577__A4 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1700_ _0030_ clknet_leaf_51_clk ram16\[1\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1631_ _0610_ _0664_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1034__I0 ram16\[1\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1562_ _0624_ _0414_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1493_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input4_I address[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0863__I3 ram16\[11\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1829_ _0159_ clknet_leaf_32_clk ram16\[10\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1752__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0839__I0 ram16\[6\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1079__S _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0993_ ram16\[0\].rb.ram1\[0\].rc.rd ram16\[0\].rb.ram1\[0\].rc.mem _0628_ _0631_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1775__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1614_ ram16\[14\].rb.ram1\[2\].rc.rd _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1545_ _0613_ _0400_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1476_ _0369_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1494__I0 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0997__A2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1410__A3 _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1174__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1798__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1330_ _0275_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1165__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1261_ _0799_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1192_ net12 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 data_in[2] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0976_ net7 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1156__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1528_ _0398_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1459_ ram16\[11\].rb.ram1\[7\].rc.mem ram16\[11\].rb.ram1\[7\].rc.rd _0358_ _0360_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1092__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0995__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1813__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1313_ ram16\[6\].rb.ram1\[7\].rc.mem _0818_ _0815_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0897__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1244_ ram16\[6\].rb.ram1\[6\].rc.mem _0770_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1175_ _0750_ _0756_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0959_ _0609_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1377__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1129__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1836__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1540__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1862_ _0192_ clknet_leaf_40_clk ram16\[12\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput10 data_in[5] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1793_ _0123_ clknet_leaf_11_clk ram16\[7\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1359__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1227_ net6 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1709__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1158_ _0704_ _0738_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1089_ _0584_ _0601_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1859__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0892__S0 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1012_ ram16\[1\].rb.ram1\[5\].rc.rd ram16\[1\].rb.ram1\[5\].rc.mem _0642_ _0644_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0875__I1 ram16\[3\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _0244_ clknet_leaf_21_clk ram16\[15\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1845_ _0175_ clknet_leaf_26_clk ram16\[11\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0883__S0 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1776_ _0106_ clknet_leaf_10_clk ram16\[6\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1681__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1291__I1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1440__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1282__I1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1630_ _0668_ _0466_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1561_ _0417_ _0421_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1492_ _0698_ _0736_ _0267_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1273__I1 ram16\[6\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ _0158_ clknet_leaf_52_clk ram16\[9\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1759_ _0089_ clknet_leaf_7_clk ram16\[5\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1264__I1 ram16\[6\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0847__S0 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0998__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0992_ _0630_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1255__I1 ram16\[6\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1069__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1613_ _0431_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1544_ _0404_ _0410_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1475_ ram16\[11\].rb.ram1\[2\].rc.mem _0786_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0997__A3 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1246__I1 ram16\[6\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1410__A4 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1260_ _0809_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1191_ _0761_ _0766_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput8 data_in[3] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1625__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1228__I1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0975_ _0619_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1892__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1463__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1527_ ram16\[12\].rb.ram1\[0\].rc.rd ram16\[12\].rb.ram1\[0\].rc.mem _0394_ _0398_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1458_ _0359_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1389_ _0313_ _0314_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1616__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1092__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1219__I1 ram16\[5\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0978__I0 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1312_ _0264_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0897__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1243_ _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1174_ ram16\[4\].rb.ram1\[4\].rc.rd _0747_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0958_ ram16\[0\].rb.ram1\[7\].rc.rd ram16\[0\].rb.ram1\[7\].rc.mem _0607_ _0609_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0889_ ram16\[0\].rb.ram1\[5\].rc.rd ram16\[1\].rb.ram1\[5\].rc.rd ram16\[8\].rb.ram1\[5\].rc.rd
+ ram16\[9\].rb.ram1\[5\].rc.rd _0546_ _0522_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1788__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1278__S _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1861_ _0191_ clknet_leaf_36_clk ram16\[12\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput11 data_in[6] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1792_ _0122_ clknet_leaf_9_clk ram16\[7\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1226_ _0789_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1157_ _0743_ _0744_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1088_ _0524_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1803__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1038__A2 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0892__S1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1349__I0 ram16\[8\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1360__I _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1011_ _0643_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1521__I0 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1913_ _0243_ clknet_leaf_18_clk ram16\[15\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0883__S1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1844_ _0174_ clknet_leaf_1_clk ram16\[10\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1775_ _0105_ clknet_leaf_10_clk ram16\[6\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1209_ _0778_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1826__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1270__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1512__I0 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1440__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1503__I0 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0857__I2 ram16\[8\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1431__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1560_ ram16\[13\].rb.ram1\[3\].rc.rd _0409_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1491_ _0377_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1355__I _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0942__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1291__S _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1849__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ _0157_ clknet_leaf_46_clk ram16\[8\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1466__S _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1758_ _0088_ clknet_leaf_13_clk ram16\[5\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0933__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1689_ _0019_ clknet_leaf_39_clk ram16\[1\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1661__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0847__S1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0924__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1652__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0991_ ram16\[0\].rb.ram1\[1\].rc.rd ram16\[0\].rb.ram1\[1\].rc.mem _0628_ _0630_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1286__S _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1612_ _0454_ _0455_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1543_ ram16\[13\].rb.ram1\[6\].rc.rd _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1474_ _0357_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1634__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1398__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1190_ ram16\[4\].rb.ram1\[1\].rc.rd _0762_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 data_in[4] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1625__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0974_ ram16\[0\].rb.ram1\[4\].rc.rd ram16\[0\].rb.ram1\[4\].rc.mem _0614_ _0619_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1526_ _0397_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1457_ ram16\[11\].rb.ram1\[6\].rc.mem _0770_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1388_ ram16\[9\].rb.ram1\[2\].rc.mem _0310_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1616__A2 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1628__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1311_ ram16\[7\].rb.ram1\[1\].rc.mem ram16\[7\].rb.ram1\[1\].rc.rd _0262_ _0264_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1363__I _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1242_ _0513_ _0501_ _0508_ _0771_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_92_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1173_ _0753_ _0755_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_44_clk clknet_2_0__leaf_clk clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0957_ _0608_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0888_ _0520_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1509_ ram16\[12\].rb.ram1\[4\].rc.rd ram16\[12\].rb.ram1\[4\].rc.mem _0384_ _0388_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0896__I0 ram16\[0\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_clk clknet_2_1__leaf_clk clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_26_clk clknet_2_3__leaf_clk clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1300__I1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1860_ _0190_ clknet_leaf_5_clk ram16\[11\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1791_ _0121_ clknet_leaf_9_clk ram16\[7\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput12 data_in[7] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1358__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_51_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1093__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1225_ ram16\[5\].rb.ram1\[3\].rc.mem ram16\[5\].rb.ram1\[3\].rc.rd _0787_ _0789_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1156_ ram16\[4\].rb.ram1\[7\].rc.mem _0741_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_17_clk clknet_2_3__leaf_clk clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1087_ net11 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1755__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_19_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0869__I0 ram16\[6\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1641__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1010_ _0641_ ram16\[1\].rb.ram1\[4\].rc.mem _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0875__I3 ram16\[11\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ _0242_ clknet_leaf_21_clk ram16\[15\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1778__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1843_ _0173_ clknet_leaf_41_clk ram16\[0\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1774_ _0104_ clknet_leaf_12_clk ram16\[6\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1208_ ram16\[5\].rb.ram1\[6\].rc.mem ram16\[5\].rb.ram1\[6\].rc.rd _0773_ _0778_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1139_ ram16\[3\].rb.ram1\[1\].rc.rd _0726_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1028__I0 ram16\[1\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1920__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1195__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1490_ ram16\[11\].rb.ram1\[0\].rc.mem ram16\[11\].rb.ram1\[0\].rc.rd _0373_ _0377_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1826_ _0156_ clknet_leaf_52_clk ram16\[9\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1757_ _0087_ clknet_leaf_7_clk ram16\[5\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1688_ _0018_ clknet_leaf_35_clk ram16\[1\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1281__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I data_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1110__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1456__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1177__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0924__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0990_ _0629_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1611_ ram16\[14\].rb.ram1\[1\].rc.mem _0448_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1542_ _0399_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1473_ _0367_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I address[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1477__S _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1809_ _0139_ clknet_leaf_51_clk ram16\[8\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1159__A2 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1403__I0 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1398__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1839__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1297__S _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0973_ _0618_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1525_ ram16\[11\].rb.ram1\[7\].rc.mem _0818_ _0373_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1456_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1387_ _0719_ _0308_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0884__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1543__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1310_ _0263_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1241_ _0798_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1172_ ram16\[4\].rb.ram1\[3\].rc.mem _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0956_ _0600_ ram16\[0\].rb.ram1\[6\].rc.mem _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0887_ _0502_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1534__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1508_ _0387_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__S _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1439_ _0343_ _0347_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1684__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0896__I1 ram16\[1\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1790_ _0120_ clknet_leaf_12_clk ram16\[7\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput13 rd_wr net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1224_ _0788_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1155_ ram16\[4\].rb.ram1\[7\].rc.rd _0738_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1086_ _0691_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0939_ ram16\[6\].rb.ram1\[0\].rc.rd ram16\[7\].rb.ram1\[0\].rc.rd ram16\[14\].rb.ram1\[0\].rc.rd
+ ram16\[15\].rb.ram1\[0\].rc.rd _0521_ _0558_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_2__f_clk clknet_0_clk clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ _0241_ clknet_leaf_20_clk ram16\[15\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1842_ _0172_ clknet_leaf_1_clk ram16\[10\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1773_ _0103_ clknet_leaf_10_clk ram16\[6\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1207_ _0777_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1138_ _0729_ _0730_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1069_ _0671_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1276__I1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1722__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0911__I _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1664__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_50_clk_I clknet_2_0__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_18_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1407__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1895__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1825_ _0155_ clknet_leaf_52_clk ram16\[9\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1756_ _0086_ clknet_leaf_25_clk ram16\[5\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1687_ _0017_ clknet_leaf_38_clk ram16\[1\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0906__I _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0999__I0 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1610_ _0624_ _0446_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1541_ _0407_ _0408_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1472_ ram16\[11\].rb.ram1\[4\].rc.mem ram16\[11\].rb.ram1\[4\].rc.rd _0363_ _0367_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1382__I _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0923__I0 ram16\[0\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1479__I1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1808_ _0138_ clknet_leaf_50_clk ram16\[8\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1739_ _0069_ clknet_leaf_3_clk ram16\[4\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1910__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0972_ _0617_ ram16\[0\].rb.ram1\[3\].rc.mem _0614_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1524_ _0396_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1455_ _0698_ _0694_ _0661_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_68_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1386_ _0306_ _0312_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1806__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1197__I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1240_ ram16\[5\].rb.ram1\[0\].rc.mem ram16\[5\].rb.ram1\[0\].rc.rd _0794_ _0798_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1171_ _0740_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0955_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0886_ _0493_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1507_ _0645_ ram16\[12\].rb.ram1\[3\].rc.mem _0384_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0895__B _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1438_ ram16\[10\].rb.ram1\[3\].rc.rd _0335_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1829__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1369_ _0704_ _0292_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0896__I2 ram16\[8\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0914__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1223_ ram16\[5\].rb.ram1\[2\].rc.mem _0786_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1154_ _0739_ _0742_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1085_ ram16\[2\].rb.ram1\[0\].rc.rd ram16\[2\].rb.ram1\[0\].rc.mem _0687_ _0691_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0938_ _0583_ _0587_ _0589_ _0591_ net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0869_ ram16\[6\].rb.ram1\[6\].rc.rd ram16\[7\].rb.ram1\[6\].rc.rd ram16\[14\].rb.ram1\[6\].rc.rd
+ ram16\[15\].rb.ram1\[6\].rc.rd _0495_ _0498_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1006__S _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1910_ _0240_ clknet_leaf_18_clk ram16\[15\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1841_ _0171_ clknet_leaf_3_clk ram16\[10\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1772_ _0102_ clknet_leaf_23_clk ram16\[6\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1674__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1206_ ram16\[5\].rb.ram1\[5\].rc.mem _0776_ _0773_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1137_ ram16\[3\].rb.ram1\[0\].rc.mem _0716_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1068_ _0681_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1496__S _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1113__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1664__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1697__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1824_ _0154_ clknet_leaf_52_clk ram16\[9\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1755_ _0085_ clknet_leaf_13_clk ram16\[5\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1686_ _0016_ clknet_leaf_42_clk ram16\[1\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0941__I1 ram16\[5\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__A2 _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0909__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1637__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1540_ ram16\[13\].rb.ram1\[5\].rc.mem _0403_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1471_ _0366_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1712__CLK clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0923__I1 ram16\[1\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1807_ _0137_ clknet_leaf_51_clk ram16\[8\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1738_ _0068_ clknet_leaf_27_clk ram16\[4\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1669_ _0300_ _0490_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1619__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1735__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1483__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1885__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0971_ net8 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1523_ ram16\[12\].rb.ram1\[1\].rc.rd ram16\[12\].rb.ram1\[1\].rc.mem _0394_ _0396_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1454_ _0353_ _0356_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1385_ ram16\[9\].rb.ram1\[4\].rc.rd _0303_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_47_clk clknet_2_0__leaf_clk clknet_leaf_47_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1085__I0 ram16\[2\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1758__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0899__I0 ram16\[2\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_38_clk clknet_2_1__leaf_clk clknet_leaf_38_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1076__I0 ram16\[2\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1170_ _0713_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_29_clk clknet_2_3__leaf_clk clknet_leaf_29_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1900__CLK clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1067__I0 ram16\[2\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0954_ _0602_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0885_ ram16\[2\].rb.ram1\[5\].rc.rd ram16\[3\].rb.ram1\[5\].rc.rd ram16\[10\].rb.ram1\[5\].rc.rd
+ ram16\[11\].rb.ram1\[5\].rc.rd _0514_ _0516_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1506_ _0386_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1437_ _0345_ _0346_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1368_ _0299_ _0300_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1299_ _0821_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1058__I0 ram16\[2\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0930__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1923__CLK clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1222_ _0772_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1153_ ram16\[4\].rb.ram1\[6\].rc.mem _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1084_ _0690_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0937_ _0555_ _0590_ _0572_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0868_ _0500_ _0511_ _0518_ _0527_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1581__I _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1451__I0 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0890__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1840_ _0170_ clknet_leaf_3_clk ram16\[10\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1771_ _0101_ clknet_leaf_12_clk ram16\[6\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1819__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1370__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1205_ net10 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1136_ _0728_ _0714_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0881__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1067_ ram16\[2\].rb.ram1\[4\].rc.rd ram16\[2\].rb.ram1\[4\].rc.mem _0677_ _0681_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1017__S _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1104__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1407__A3 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1823_ _0153_ clknet_leaf_52_clk ram16\[9\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1791__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1754_ _0084_ clknet_leaf_25_clk ram16\[5\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1040__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1591__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1685_ _0015_ clknet_leaf_35_clk ram16\[1\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0941__I2 ram16\[12\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1119_ _0715_ _0717_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1300__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1582__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0932__I2 ram16\[12\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1098__A1 ram16\[3\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1470_ ram16\[11\].rb.ram1\[3\].rc.mem _0783_ _0363_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0923__I2 ram16\[8\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1089__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1806_ _0136_ clknet_leaf_48_clk ram16\[8\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1737_ _0067_ clknet_leaf_32_clk ram16\[4\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1668_ _0659_ _0318_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1599_ _0617_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1555__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0843__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0970_ _0616_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1546__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0395_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1453_ ram16\[10\].rb.ram1\[0\].rc.rd _0350_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1384_ _0309_ _0311_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1537__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0899__I1 ram16\[3\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1702__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1852__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0838__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0953_ _0505_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_0884_ _0503_ _0541_ _0510_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1505_ ram16\[12\].rb.ram1\[5\].rc.rd ram16\[12\].rb.ram1\[5\].rc.mem _0384_ _0386_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1436_ ram16\[10\].rb.ram1\[2\].rc.mem _0342_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1367_ ram16\[9\].rb.ram1\[7\].rc.mem _0297_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1298_ _0256_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1455__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0889__S0 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_2_0__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_16_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1446__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1221_ net7 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1748__CLK clknet_leaf_6_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1152_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1083_ _0659_ ram16\[1\].rb.ram1\[7\].rc.mem _0656_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1898__CLK clknet_leaf_20_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0936_ ram16\[2\].rb.ram1\[1\].rc.rd ram16\[3\].rb.ram1\[1\].rc.rd ram16\[10\].rb.ram1\[1\].rc.rd
+ ram16\[11\].rb.ram1\[1\].rc.rd _0504_ _0570_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0867_ _0519_ _0523_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1212__I1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1419_ _0333_ _0334_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1203__I1 ram16\[5\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1667__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1770_ _0100_ clknet_leaf_23_clk ram16\[6\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1204_ _0775_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1135_ net5 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0881__A2 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1066_ _0680_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1899_ _0229_ clknet_leaf_12_clk ram16\[14\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0919_ ram16\[6\].rb.ram1\[2\].rc.rd ram16\[7\].rb.ram1\[2\].rc.rd ram16\[14\].rb.ram1\[2\].rc.rd
+ ram16\[15\].rb.ram1\[2\].rc.rd _0537_ _0558_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__1913__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1208__S _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0846__I _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1822_ _0152_ clknet_leaf_44_clk ram16\[9\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1753_ _0083_ clknet_leaf_25_clk ram16\[5\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1684_ _0014_ clknet_leaf_0_clk ram16\[0\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1118_ ram16\[3\].rb.ram1\[3\].rc.mem _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1049_ _0584_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_41_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1028__S _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1809__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1342__I0 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1098__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1333__I0 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1200__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1805_ _0135_ clknet_leaf_50_clk ram16\[8\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1736_ _0066_ clknet_leaf_27_clk ram16\[4\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1667_ _0486_ _0489_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1598_ _0431_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1311__S _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1020__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1521_ _0655_ ram16\[12\].rb.ram1\[0\].rc.mem _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1452_ _0355_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1383_ ram16\[9\].rb.ram1\[3\].rc.mem _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1719_ _0049_ clknet_leaf_33_clk ram16\[3\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1306__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1105__I _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0854__I _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0952_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_0883_ ram16\[4\].rb.ram1\[5\].rc.rd ram16\[5\].rb.ram1\[5\].rc.rd ram16\[12\].rb.ram1\[5\].rc.rd
+ ram16\[13\].rb.ram1\[5\].rc.rd _0540_ _0506_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1504_ _0385_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1527__I0 ram16\[12\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1435_ _0719_ _0340_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1366_ ram16\[9\].rb.ram1\[7\].rc.rd _0292_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1297_ ram16\[7\].rb.ram1\[4\].rc.mem ram16\[7\].rb.ram1\[4\].rc.rd _0827_ _0256_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1455__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0889__S1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1518__I0 ram16\[12\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1446__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0849__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1509__I0 ram16\[12\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1220_ _0785_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1151_ _0735_ _0525_ _0603_ _0736_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1082_ _0689_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0935_ _0545_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0866_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1418_ ram16\[10\].rb.ram1\[5\].rc.mem _0329_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1349_ ram16\[8\].rb.ram1\[1\].rc.rd ram16\[8\].rb.ram1\[1\].rc.mem _0284_ _0286_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1842__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1715__CLK clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1203_ ram16\[5\].rb.ram1\[7\].rc.mem ram16\[5\].rb.ram1\[7\].rc.rd _0773_ _0775_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_15_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1134_ _0721_ _0727_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1065_ _0645_ ram16\[2\].rb.ram1\[3\].rc.mem _0677_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1898_ _0228_ clknet_leaf_20_clk ram16\[14\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0918_ _0560_ _0565_ _0569_ _0573_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_0849_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1649__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0880__I0 ram16\[6\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1888__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0943__S0 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0862__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1821_ _0151_ clknet_leaf_52_clk ram16\[9\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1752_ _0082_ clknet_leaf_26_clk ram16\[5\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1683_ _0013_ clknet_leaf_0_clk ram16\[0\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1351__I1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0934__S0 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1117_ _0699_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1048_ _0669_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1309__S _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1108__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0925__S0 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1219__S _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1903__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1804_ _0134_ clknet_leaf_40_clk ram16\[8\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1735_ _0065_ clknet_leaf_32_clk ram16\[4\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ ram16\[15\].rb.ram1\[0\].rc.rd _0480_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1597_ _0440_ _0445_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1021__I0 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0907__S0 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1324__I1 ram16\[8\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1598__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1012__I0 ram16\[1\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1079__I0 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1520_ _0378_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1451_ _0732_ ram16\[0\].rb.ram1\[7\].rc.mem _0628_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1382_ _0296_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1306__I1 ram16\[7\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1211__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1718_ _0048_ clknet_leaf_43_clk ram16\[3\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1649_ ram16\[15\].rb.ram1\[2\].rc.mem _0475_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0899__I3 ram16\[11\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1170__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1322__S _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0960__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1031__I _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0951_ net13 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0882_ _0494_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1503_ _0641_ ram16\[12\].rb.ram1\[4\].rc.mem _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1434_ _0338_ _0344_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1365_ _0293_ _0298_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1296_ _0830_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1142__S _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1455__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1771__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0955__I _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1052__S _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1150_ _0692_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0893__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1081_ ram16\[2\].rb.ram1\[1\].rc.rd ram16\[2\].rb.ram1\[1\].rc.mem _0687_ _0689_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1794__CLK clknet_leaf_10_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0934_ ram16\[0\].rb.ram1\[1\].rc.rd ram16\[1\].rb.ram1\[1\].rc.rd ram16\[8\].rb.ram1\[1\].rc.rd
+ ram16\[9\].rb.ram1\[1\].rc.rd _0566_ _0567_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0865_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1373__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1417_ _0704_ _0326_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1348_ _0285_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1279_ _0820_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1047__S _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1364__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1116__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1202_ _0774_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1133_ ram16\[3\].rb.ram1\[2\].rc.rd _0726_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1064_ _0679_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1043__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0917_ _0545_ _0571_ _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1594__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1897_ _0227_ clknet_leaf_20_clk ram16\[14\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0848_ net3 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1585__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1505__S _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0943__S1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1240__S _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0871__I1 ram16\[5\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1820_ _0150_ clknet_leaf_43_clk ram16\[9\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1751_ _0081_ clknet_leaf_24_clk ram16\[5\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1682_ _0012_ clknet_leaf_0_clk ram16\[0\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1832__CLK clknet_leaf_32_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1116_ _0713_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0934__S1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1047_ ram16\[1\].rb.ram1\[0\].rc.rd ram16\[1\].rb.ram1\[0\].rc.mem _0656_ _0669_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_14_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1855__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1558__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1803_ _0133_ clknet_leaf_47_clk ram16\[8\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1734_ _0064_ clknet_leaf_30_clk ram16\[4\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1665_ _0438_ _0488_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1596_ ram16\[14\].rb.ram1\[5\].rc.rd _0441_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0907__S1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1450_ _0349_ _0354_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1381_ _0713_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1717_ _0047_ clknet_leaf_33_clk ram16\[3\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1648_ _0620_ _0473_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1579_ _0600_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1481__I1 ram16\[11\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0950_ _0520_ _0601_ _0524_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1621__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1472__I1 ram16\[11\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0881_ _0536_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1502_ _0378_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1433_ ram16\[10\].rb.ram1\[4\].rc.rd _0335_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0983__I0 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1364_ ram16\[9\].rb.ram1\[6\].rc.mem _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1295_ ram16\[7\].rb.ram1\[3\].rc.mem _0783_ _0827_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1222__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1463__I1 ram16\[11\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1916__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0974__I0 ram16\[0\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1333__S _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1132__I _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0971__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1206__I1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0893__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1080_ _0688_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1142__I0 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0933_ _0561_ _0586_ _0564_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_0864_ net3 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0956__I0 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1416_ _0331_ _0332_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1347_ _0655_ ram16\[8\].rb.ram1\[0\].rc.mem _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1278_ ram16\[6\].rb.ram1\[0\].rc.mem ram16\[6\].rb.ram1\[0\].rc.rd _0815_ _0820_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0966__I _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1063__S _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1201_ ram16\[5\].rb.ram1\[6\].rc.mem _0770_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1132_ _0695_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1063_ ram16\[2\].rb.ram1\[5\].rc.rd ram16\[2\].rb.ram1\[5\].rc.mem _0677_ _0679_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1761__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1043__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0916_ _0525_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1896_ _0226_ clknet_leaf_20_clk ram16\[14\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0847_ ram16\[4\].rb.ram1\[7\].rc.rd ram16\[5\].rb.ram1\[7\].rc.rd ram16\[12\].rb.ram1\[7\].rc.rd
+ ram16\[13\].rb.ram1\[7\].rc.rd _0504_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1058__S _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1521__S _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1750_ _0080_ clknet_leaf_17_clk ram16\[5\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__0871__I2 ram16\[12\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1681_ _0011_ clknet_leaf_0_clk ram16\[0\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input9_I data_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1115_ _0695_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1046_ _0665_ _0668_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1879_ _0209_ clknet_leaf_29_clk ram16\[13\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1516__S _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_3__f_clk clknet_0_clk clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1802_ _0132_ clknet_leaf_42_clk ram16\[8\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1733_ _0063_ clknet_leaf_32_clk ram16\[4\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1664_ _0659_ _0456_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1595_ _0443_ _0444_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1029_ _0654_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_2_3__f_clk_I clknet_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1135__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0920__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1822__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1246__S _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1380_ _0291_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1716_ _0046_ clknet_leaf_48_clk ram16\[2\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1647_ _0471_ _0477_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1578_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1845__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_28_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1449__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1621__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0880_ ram16\[6\].rb.ram1\[5\].rc.rd ram16\[7\].rb.ram1\[5\].rc.rd ram16\[14\].rb.ram1\[5\].rc.rd
+ ram16\[15\].rb.ram1\[5\].rc.rd _0537_ _0498_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__1718__CLK clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0879__I _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1501_ _0383_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1432_ _0341_ _0343_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1868__CLK clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1363_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1294_ _0829_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1603__A2 _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0932_ ram16\[4\].rb.ram1\[1\].rc.rd ram16\[5\].rb.ram1\[1\].rc.rd ram16\[12\].rb.ram1\[1\].rc.rd
+ ram16\[13\].rb.ram1\[1\].rc.rd _0585_ _0562_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_clk clknet_2_1__leaf_clk clknet_leaf_40_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0863_ ram16\[2\].rb.ram1\[7\].rc.rd ram16\[3\].rb.ram1\[7\].rc.rd ram16\[10\].rb.ram1\[7\].rc.rd
+ ram16\[11\].rb.ram1\[7\].rc.rd _0521_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1690__CLK clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1415_ ram16\[10\].rb.ram1\[7\].rc.mem _0329_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1346_ _0268_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_84_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1277_ _0819_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1233__I _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_31_clk clknet_2_1__leaf_clk clknet_leaf_31_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1408__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1344__S _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0982__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk clknet_leaf_22_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1200_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1131_ _0724_ _0725_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1906__CLK clknet_leaf_9_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1062_ _0678_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1579__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk clknet_leaf_13_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_0915_ ram16\[0\].rb.ram1\[3\].rc.rd ram16\[1\].rb.ram1\[3\].rc.rd ram16\[8\].rb.ram1\[3\].rc.rd
+ ram16\[9\].rb.ram1\[3\].rc.rd _0546_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1895_ _0225_ clknet_leaf_19_clk ram16\[14\].rb.ram1\[5\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0846_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1329_ _0641_ ram16\[8\].rb.ram1\[4\].rc.mem _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0977__I _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1074__S _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0928__S0 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ _0010_ clknet_leaf_0_clk ram16\[0\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0887__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0919__S0 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk clknet_leaf_2_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1114_ net8 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1045_ ram16\[15\].rb.ram1\[7\].rc.mem _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1511__I _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1878_ _0208_ clknet_leaf_16_clk ram16\[13\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1015__I0 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1801_ _0131_ clknet_leaf_40_clk ram16\[8\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1732_ _0062_ clknet_leaf_2_clk ram16\[3\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ _0483_ _0487_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1006__I0 ram16\[1\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1594_ ram16\[14\].rb.ram1\[4\].rc.mem _0435_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1182__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1309__I1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1028_ ram16\[1\].rb.ram1\[2\].rc.rd ram16\[1\].rb.ram1\[2\].rc.mem _0649_ _0654_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1774__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0920__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1527__S _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1164__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1262__S _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1797__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1715_ _0045_ clknet_leaf_46_clk ram16\[1\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1646_ ram16\[15\].rb.ram1\[4\].rc.rd _0465_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1577_ _0585_ _0294_ _0633_ _0661_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1155__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1347__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1146__I _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1257__S _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1385__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ ram16\[12\].rb.ram1\[6\].rc.rd ram16\[12\].rb.ram1\[6\].rc.mem _0379_ _0383_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1431_ ram16\[10\].rb.ram1\[3\].rc.mem _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1137__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1362_ _0495_ _0294_ _0509_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1293_ ram16\[7\].rb.ram1\[5\].rc.mem ram16\[7\].rb.ram1\[5\].rc.rd _0827_ _0829_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1376__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ ram16\[15\].rb.ram1\[7\].rc.rd _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1812__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1367__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0931_ _0584_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_12_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0862_ _0497_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1835__CLK clknet_leaf_3_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_27_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1414_ ram16\[10\].rb.ram1\[7\].rc.rd _0326_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1345_ _0283_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1276_ ram16\[5\].rb.ram1\[7\].rc.mem _0818_ _0794_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1708__CLK clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0883__I1 ram16\[5\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1037__A1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1588__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__CLK clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1130_ ram16\[3\].rb.ram1\[1\].rc.mem _0716_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1061_ _0641_ ram16\[2\].rb.ram1\[4\].rc.mem _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1579__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1894_ _0224_ clknet_leaf_18_clk ram16\[14\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0914_ _0497_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0845_ net4 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1328_ _0268_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1259_ ram16\[6\].rb.ram1\[4\].rc.mem ram16\[6\].rb.ram1\[4\].rc.rd _0805_ _0809_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0873__S0 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0928__S1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1680__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0942__B _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0919__S1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1113_ _0706_ _0712_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1044_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0847__I1 ram16\[5\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1877_ _0207_ clknet_leaf_29_clk ram16\[13\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1488__A1 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0988__I _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1085__S _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1800_ _0130_ clknet_leaf_35_clk ram16\[8\].rb.ram1\[6\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1731_ _0061_ clknet_leaf_41_clk ram16\[2\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1662_ ram16\[15\].rb.ram1\[1\].rc.rd _0480_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1593_ _0613_ _0432_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1027_ _0653_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1642__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1919__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1484__I1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1475__I1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1714_ _0044_ clknet_leaf_48_clk ram16\[2\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1645_ _0474_ _0476_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1576_ _0427_ _0430_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1252__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1741__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1466__I1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1891__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1457__I1 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1337__I _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ _0328_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1361_ _0267_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1273__S _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1292_ _0828_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1764__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1628_ _0663_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1559_ _0419_ _0420_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0996__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1787__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0930_ net1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1268__S _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0861_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1413_ _0327_ _0330_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1344_ ram16\[8\].rb.ram1\[2\].rc.rd ram16\[8\].rb.ram1\[2\].rc.mem _0279_ _0283_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1275_ net12 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0883__I2 ram16\[12\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1060_ _0671_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1893_ _0223_ clknet_leaf_18_clk ram16\[14\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0913_ _0493_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_0844_ _0494_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1461__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1327_ _0273_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1258_ _0808_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1189_ _0764_ _0765_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0873__S1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0950__A1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_11_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1825__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1112_ ram16\[3\].rb.ram1\[5\].rc.rd _0707_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1043_ _0660_ _0661_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0847__I2 ram16\[12\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1876_ _0206_ clknet_leaf_51_clk ram16\[12\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1421__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1848__CLK clknet_leaf_26_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1488__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1660__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1412__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1176__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ _0060_ clknet_leaf_2_clk ram16\[3\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1661_ _0485_ _0486_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1276__S _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1592_ _0436_ _0442_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I data_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1026_ _0652_ ram16\[1\].rb.ram1\[1\].rc.mem _0649_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1642__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1859_ _0189_ clknet_leaf_43_clk ram16\[10\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1158__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1713_ _0043_ clknet_leaf_48_clk ram16\[2\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1693__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1644_ ram16\[15\].rb.ram1\[3\].rc.mem _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1575_ ram16\[13\].rb.ram1\[0\].rc.rd _0424_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1009_ _0634_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1551__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1443__I _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1606__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_52_clk clknet_2_0__leaf_clk clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1360_ _0501_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1291_ ram16\[7\].rb.ram1\[4\].rc.mem _0779_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1909__CLK clknet_leaf_17_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_43_clk clknet_2_1__leaf_clk clknet_leaf_43_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1081__I0 ram16\[2\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _0463_ _0464_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1558_ ram16\[13\].rb.ram1\[2\].rc.mem _0416_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1489_ _0332_ _0376_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_34_clk clknet_2_1__leaf_clk clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1072__I0 ram16\[2\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0860_ net1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1063__I0 ram16\[2\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1284__S _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1412_ ram16\[10\].rb.ram1\[6\].rc.mem _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1731__CLK clknet_leaf_41_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1343_ _0282_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1274_ _0817_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_16_clk clknet_2_3__leaf_clk clknet_leaf_16_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1459__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0989_ _0627_ ram16\[0\].rb.ram1\[0\].rc.mem _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1054__I0 ram16\[2\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1754__CLK clknet_leaf_25_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _0222_ clknet_leaf_6_clk ram16\[13\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0912_ ram16\[2\].rb.ram1\[3\].rc.rd ram16\[3\].rb.ram1\[3\].rc.rd ram16\[10\].rb.ram1\[3\].rc.rd
+ ram16\[11\].rb.ram1\[3\].rc.rd _0566_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_0843_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1078__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk clknet_leaf_5_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1326_ ram16\[8\].rb.ram1\[6\].rc.rd ram16\[8\].rb.ram1\[6\].rc.mem _0269_ _0273_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1257_ ram16\[6\].rb.ram1\[3\].rc.mem _0783_ _0805_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1188_ ram16\[4\].rb.ram1\[0\].rc.mem _0754_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1777__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1111_ _0710_ _0711_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1042_ _0659_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1875_ _0205_ clknet_leaf_16_clk ram16\[11\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1185__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1472__S _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1309_ ram16\[7\].rb.ram1\[0\].rc.mem _0793_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1496__I0 ram16\[12\].rb.ram1\[7\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1176__A2 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ ram16\[15\].rb.ram1\[0\].rc.mem _0475_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1591_ ram16\[14\].rb.ram1\[6\].rc.rd _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1167__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1091__I _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1025_ net6 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_10_clk_I clknet_2_2__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1858_ _0188_ clknet_leaf_5_clk ram16\[11\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1789_ _0119_ clknet_leaf_9_clk ram16\[7\].rb.ram1\[2\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1815__CLK clknet_leaf_34_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1158__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_25_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1094__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1838__CLK clknet_leaf_44_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1712_ _0042_ clknet_leaf_47_clk ram16\[2\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1388__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1643_ _0666_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _0429_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1560__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1008_ net9 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1551__A2 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1290_ _0821_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1626_ ram16\[15\].rb.ram1\[6\].rc.mem _0667_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1557_ _0620_ _0414_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1488_ _0767_ _0350_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1683__CLK clknet_leaf_0_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0894__S0 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1411_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1342_ _0652_ ram16\[8\].rb.ram1\[1\].rc.mem _0279_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1273_ ram16\[6\].rb.ram1\[1\].rc.mem ram16\[6\].rb.ram1\[1\].rc.rd _0815_ _0817_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0885__S0 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0988_ _0606_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1475__S _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1609_ _0449_ _0453_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ _0221_ clknet_leaf_41_clk ram16\[12\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_0911_ _0515_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0842_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1295__S _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1325_ _0272_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1256_ _0807_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1187_ _0728_ _0752_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1721__CLK clknet_leaf_33_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1266__I1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1871__CLK clknet_leaf_51_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1110_ ram16\[3\].rb.ram1\[4\].rc.mem _0700_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1041_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1257__I1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1874_ _0204_ clknet_leaf_51_clk ram16\[12\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1308_ _0821_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1239_ _0744_ _0797_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1744__CLK clknet_leaf_1_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1248__I1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1894__CLK clknet_leaf_18_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1636__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1590_ _0431_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1573__S _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1372__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1024_ _0651_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0989__I0 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1857_ _0187_ clknet_leaf_5_clk ram16\[11\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1788_ _0118_ clknet_leaf_20_clk ram16\[7\].rb.ram1\[4\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1094__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1192__I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1711_ _0041_ clknet_leaf_48_clk ram16\[2\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1642_ _0617_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1573_ _0732_ ram16\[12\].rb.ram1\[7\].rc.mem _0394_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1007_ _0640_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1320__I0 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1909_ _0239_ clknet_leaf_17_clk ram16\[15\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1805__CLK clknet_leaf_50_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_24_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_39_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1625_ _0600_ _0664_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1556_ _0412_ _0418_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1487_ _0375_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1001__S _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1828__CLK clknet_leaf_52_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0894__S1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1410_ _0289_ _0290_ _0509_ _0295_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1341_ _0281_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1272_ _0816_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1380__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1523__I0 ram16\[12\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0885__S1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0987_ net5 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1608_ ram16\[14\].rb.ram1\[3\].rc.rd _0441_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1539_ _0610_ _0400_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1290__I _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1514__I0 ram16\[12\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1465__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0953__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1505__I0 ram16\[12\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0910_ _0513_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1890_ _0220_ clknet_leaf_6_clk ram16\[13\].rb.ram1\[1\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1433__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0841_ net2 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XANTENNA__0944__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1324_ _0638_ ram16\[8\].rb.ram1\[5\].rc.mem _0269_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1255_ ram16\[6\].rb.ram1\[5\].rc.mem ram16\[6\].rb.ram1\[5\].rc.rd _0805_ _0807_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1186_ _0758_ _0763_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1424__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1486__S _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0935__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1673__CLK clknet_leaf_39_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1415__A2 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0926__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1040_ _0660_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__A2 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1873_ _0203_ clknet_leaf_51_clk ram16\[12\].rb.ram1\[0\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1696__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0917__A1 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1307_ _0261_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1238_ _0767_ _0762_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1169_ _0737_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1636__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1023_ ram16\[1\].rb.ram1\[3\].rc.rd ram16\[1\].rb.ram1\[3\].rc.mem _0649_ _0651_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1925_ _0255_ clknet_leaf_44_clk ram16\[9\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1856_ _0186_ clknet_leaf_14_clk ram16\[11\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1787_ _0117_ clknet_leaf_12_clk ram16\[7\].rb.ram1\[3\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1711__CLK clknet_leaf_48_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input13_I rd_wr vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1004__S _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0921__S0 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0912__S0 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1710_ _0040_ clknet_leaf_47_clk ram16\[2\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1641_ _0663_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1545__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1572_ _0423_ _0428_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1734__CLK clknet_leaf_30_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I data_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_46_clk clknet_2_0__leaf_clk clknet_leaf_46_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1006_ ram16\[1\].rb.ram1\[6\].rc.rd ram16\[1\].rb.ram1\[6\].rc.mem _0635_ _0640_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0903__S0 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1320__I1 ram16\[8\].rb.ram1\[6\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1908_ _0238_ clknet_leaf_9_clk ram16\[14\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1839_ _0169_ clknet_leaf_1_clk ram16\[10\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1494__S _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1757__CLK clknet_leaf_7_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_28_clk clknet_2_3__leaf_clk clknet_leaf_28_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1624_ _0459_ _0462_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1555_ ram16\[13\].rb.ram1\[4\].rc.rd _0409_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1486_ ram16\[11\].rb.ram1\[1\].rc.mem ram16\[11\].rb.ram1\[1\].rc.rd _0373_ _0375_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk clknet_leaf_19_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1340_ ram16\[8\].rb.ram1\[3\].rc.rd ram16\[8\].rb.ram1\[3\].rc.mem _0279_ _0281_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1271_ ram16\[6\].rb.ram1\[0\].rc.mem _0793_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1922__CLK clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0986_ _0626_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk clknet_leaf_8_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_1607_ _0451_ _0452_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1538_ _0405_ _0406_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1469_ _0365_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1012__S _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_23_clk_I clknet_2_3__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1130__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_clk_I clknet_2_1__leaf_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0840_ _0493_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__0944__A2 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1323_ _0271_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1254_ _0806_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1185_ ram16\[4\].rb.ram1\[2\].rc.rd _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0969_ ram16\[0\].rb.ram1\[5\].rc.rd ram16\[0\].rb.ram1\[5\].rc.mem _0614_ _0616_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1188__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0935__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1112__A2 _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1179__A2 _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1103__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1872_ _0202_ clknet_leaf_50_clk ram16\[12\].rb.ram1\[2\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1306_ ram16\[7\].rb.ram1\[2\].rc.mem ram16\[7\].rb.ram1\[2\].rc.rd _0257_ _0261_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1237_ _0796_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1168_ _0746_ _0751_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1099_ ram16\[3\].rb.ram1\[7\].rc.mem _0700_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1790__CLK clknet_leaf_12_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1022_ _0650_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1924_ _0254_ clknet_leaf_8_clk ram16\[15\].rb.ram1\[0\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1855_ _0185_ clknet_leaf_5_clk ram16\[11\].rb.ram1\[1\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1786_ _0116_ clknet_leaf_21_clk ram16\[7\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1563__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1094__A4 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0921__S1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0912__S1 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1242__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1640_ _0468_ _0472_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1571_ ram16\[13\].rb.ram1\[1\].rc.rd _0424_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1005_ _0639_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0903__S1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1907_ _0237_ clknet_leaf_16_clk ram16\[13\].rb.ram1\[7\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1838_ _0168_ clknet_leaf_44_clk ram16\[10\].rb.ram1\[3\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1769_ _0099_ clknet_leaf_22_clk ram16\[6\].rb.ram1\[4\].rc.mem vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1015__S _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0889__I1 ram16\[1\].rb.ram1\[5\].rc.rd vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1701__CLK clknet_leaf_35_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1623_ ram16\[14\].rb.ram1\[0\].rc.rd _0456_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1554_ _0415_ _0417_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1485_ _0374_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

