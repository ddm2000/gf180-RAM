magic
tech gf180mcuC
magscale 1 10
timestamp 1670244893
<< metal1 >>
rect 43698 96574 43710 96626
rect 43762 96623 43774 96626
rect 45042 96623 45054 96626
rect 43762 96577 45054 96623
rect 43762 96574 43774 96577
rect 45042 96574 45054 96577
rect 45106 96574 45118 96626
rect 56130 96574 56142 96626
rect 56194 96623 56206 96626
rect 56802 96623 56814 96626
rect 56194 96577 56814 96623
rect 56194 96574 56206 96577
rect 56802 96574 56814 96577
rect 56866 96574 56878 96626
rect 1344 96458 98560 96492
rect 1344 96406 4478 96458
rect 4530 96406 4582 96458
rect 4634 96406 4686 96458
rect 4738 96406 35198 96458
rect 35250 96406 35302 96458
rect 35354 96406 35406 96458
rect 35458 96406 65918 96458
rect 65970 96406 66022 96458
rect 66074 96406 66126 96458
rect 66178 96406 96638 96458
rect 96690 96406 96742 96458
rect 96794 96406 96846 96458
rect 96898 96406 98560 96458
rect 1344 96372 98560 96406
rect 6738 96126 6750 96178
rect 6802 96126 6814 96178
rect 19170 96126 19182 96178
rect 19234 96126 19246 96178
rect 31266 96126 31278 96178
rect 31330 96126 31342 96178
rect 45042 96126 45054 96178
rect 45106 96126 45118 96178
rect 56802 96126 56814 96178
rect 56866 96126 56878 96178
rect 68898 96126 68910 96178
rect 68962 96126 68974 96178
rect 81330 96126 81342 96178
rect 81394 96126 81406 96178
rect 94322 96126 94334 96178
rect 94386 96126 94398 96178
rect 8318 96066 8370 96078
rect 58382 96066 58434 96078
rect 93102 96066 93154 96078
rect 7858 96014 7870 96066
rect 7922 96014 7934 96066
rect 20290 96014 20302 96066
rect 20354 96014 20366 96066
rect 32162 96014 32174 96066
rect 32226 96014 32238 96066
rect 45938 96014 45950 96066
rect 46002 96014 46014 96066
rect 57698 96014 57710 96066
rect 57762 96014 57774 96066
rect 70018 96014 70030 96066
rect 70082 96014 70094 96066
rect 82338 96014 82350 96066
rect 82402 96014 82414 96066
rect 93874 96014 93886 96066
rect 93938 96014 93950 96066
rect 8318 96002 8370 96014
rect 58382 96002 58434 96014
rect 93102 96002 93154 96014
rect 21310 95842 21362 95854
rect 21310 95778 21362 95790
rect 33070 95842 33122 95854
rect 33070 95778 33122 95790
rect 46622 95842 46674 95854
rect 46622 95778 46674 95790
rect 70478 95842 70530 95854
rect 70478 95778 70530 95790
rect 82910 95842 82962 95854
rect 82910 95778 82962 95790
rect 1344 95674 98560 95708
rect 1344 95622 19838 95674
rect 19890 95622 19942 95674
rect 19994 95622 20046 95674
rect 20098 95622 50558 95674
rect 50610 95622 50662 95674
rect 50714 95622 50766 95674
rect 50818 95622 81278 95674
rect 81330 95622 81382 95674
rect 81434 95622 81486 95674
rect 81538 95622 98560 95674
rect 1344 95588 98560 95622
rect 1344 94890 98560 94924
rect 1344 94838 4478 94890
rect 4530 94838 4582 94890
rect 4634 94838 4686 94890
rect 4738 94838 35198 94890
rect 35250 94838 35302 94890
rect 35354 94838 35406 94890
rect 35458 94838 65918 94890
rect 65970 94838 66022 94890
rect 66074 94838 66126 94890
rect 66178 94838 96638 94890
rect 96690 94838 96742 94890
rect 96794 94838 96846 94890
rect 96898 94838 98560 94890
rect 1344 94804 98560 94838
rect 1344 94106 98560 94140
rect 1344 94054 19838 94106
rect 19890 94054 19942 94106
rect 19994 94054 20046 94106
rect 20098 94054 50558 94106
rect 50610 94054 50662 94106
rect 50714 94054 50766 94106
rect 50818 94054 81278 94106
rect 81330 94054 81382 94106
rect 81434 94054 81486 94106
rect 81538 94054 98560 94106
rect 1344 94020 98560 94054
rect 1344 93322 98560 93356
rect 1344 93270 4478 93322
rect 4530 93270 4582 93322
rect 4634 93270 4686 93322
rect 4738 93270 35198 93322
rect 35250 93270 35302 93322
rect 35354 93270 35406 93322
rect 35458 93270 65918 93322
rect 65970 93270 66022 93322
rect 66074 93270 66126 93322
rect 66178 93270 96638 93322
rect 96690 93270 96742 93322
rect 96794 93270 96846 93322
rect 96898 93270 98560 93322
rect 1344 93236 98560 93270
rect 1344 92538 98560 92572
rect 1344 92486 19838 92538
rect 19890 92486 19942 92538
rect 19994 92486 20046 92538
rect 20098 92486 50558 92538
rect 50610 92486 50662 92538
rect 50714 92486 50766 92538
rect 50818 92486 81278 92538
rect 81330 92486 81382 92538
rect 81434 92486 81486 92538
rect 81538 92486 98560 92538
rect 1344 92452 98560 92486
rect 1344 91754 98560 91788
rect 1344 91702 4478 91754
rect 4530 91702 4582 91754
rect 4634 91702 4686 91754
rect 4738 91702 35198 91754
rect 35250 91702 35302 91754
rect 35354 91702 35406 91754
rect 35458 91702 65918 91754
rect 65970 91702 66022 91754
rect 66074 91702 66126 91754
rect 66178 91702 96638 91754
rect 96690 91702 96742 91754
rect 96794 91702 96846 91754
rect 96898 91702 98560 91754
rect 1344 91668 98560 91702
rect 1344 90970 98560 91004
rect 1344 90918 19838 90970
rect 19890 90918 19942 90970
rect 19994 90918 20046 90970
rect 20098 90918 50558 90970
rect 50610 90918 50662 90970
rect 50714 90918 50766 90970
rect 50818 90918 81278 90970
rect 81330 90918 81382 90970
rect 81434 90918 81486 90970
rect 81538 90918 98560 90970
rect 1344 90884 98560 90918
rect 1344 90186 98560 90220
rect 1344 90134 4478 90186
rect 4530 90134 4582 90186
rect 4634 90134 4686 90186
rect 4738 90134 35198 90186
rect 35250 90134 35302 90186
rect 35354 90134 35406 90186
rect 35458 90134 65918 90186
rect 65970 90134 66022 90186
rect 66074 90134 66126 90186
rect 66178 90134 96638 90186
rect 96690 90134 96742 90186
rect 96794 90134 96846 90186
rect 96898 90134 98560 90186
rect 1344 90100 98560 90134
rect 1344 89402 98560 89436
rect 1344 89350 19838 89402
rect 19890 89350 19942 89402
rect 19994 89350 20046 89402
rect 20098 89350 50558 89402
rect 50610 89350 50662 89402
rect 50714 89350 50766 89402
rect 50818 89350 81278 89402
rect 81330 89350 81382 89402
rect 81434 89350 81486 89402
rect 81538 89350 98560 89402
rect 1344 89316 98560 89350
rect 68226 88958 68238 89010
rect 68290 88958 68302 89010
rect 90850 88958 90862 89010
rect 90914 88958 90926 89010
rect 63086 88898 63138 88910
rect 63086 88834 63138 88846
rect 63534 88898 63586 88910
rect 71598 88898 71650 88910
rect 68898 88846 68910 88898
rect 68962 88846 68974 88898
rect 71026 88846 71038 88898
rect 71090 88846 71102 88898
rect 91634 88846 91646 88898
rect 91698 88846 91710 88898
rect 93762 88846 93774 88898
rect 93826 88846 93838 88898
rect 63534 88834 63586 88846
rect 71598 88834 71650 88846
rect 1344 88618 98560 88652
rect 1344 88566 4478 88618
rect 4530 88566 4582 88618
rect 4634 88566 4686 88618
rect 4738 88566 35198 88618
rect 35250 88566 35302 88618
rect 35354 88566 35406 88618
rect 35458 88566 65918 88618
rect 65970 88566 66022 88618
rect 66074 88566 66126 88618
rect 66178 88566 96638 88618
rect 96690 88566 96742 88618
rect 96794 88566 96846 88618
rect 96898 88566 98560 88618
rect 1344 88532 98560 88566
rect 3266 88286 3278 88338
rect 3330 88286 3342 88338
rect 61854 88226 61906 88238
rect 62514 88174 62526 88226
rect 62578 88174 62590 88226
rect 61854 88162 61906 88174
rect 57710 88114 57762 88126
rect 63534 88114 63586 88126
rect 1922 88062 1934 88114
rect 1986 88062 1998 88114
rect 62626 88062 62638 88114
rect 62690 88062 62702 88114
rect 57710 88050 57762 88062
rect 63534 88050 63586 88062
rect 54798 88002 54850 88014
rect 54798 87938 54850 87950
rect 57374 88002 57426 88014
rect 57374 87938 57426 87950
rect 59614 88002 59666 88014
rect 59614 87938 59666 87950
rect 60622 88002 60674 88014
rect 60622 87938 60674 87950
rect 61518 88002 61570 88014
rect 61518 87938 61570 87950
rect 63870 88002 63922 88014
rect 63870 87938 63922 87950
rect 64430 88002 64482 88014
rect 64430 87938 64482 87950
rect 70478 88002 70530 88014
rect 70478 87938 70530 87950
rect 71038 88002 71090 88014
rect 71038 87938 71090 87950
rect 1344 87834 98560 87868
rect 1344 87782 19838 87834
rect 19890 87782 19942 87834
rect 19994 87782 20046 87834
rect 20098 87782 50558 87834
rect 50610 87782 50662 87834
rect 50714 87782 50766 87834
rect 50818 87782 81278 87834
rect 81330 87782 81382 87834
rect 81434 87782 81486 87834
rect 81538 87782 98560 87834
rect 1344 87748 98560 87782
rect 58046 87666 58098 87678
rect 58046 87602 58098 87614
rect 87278 87554 87330 87566
rect 54338 87502 54350 87554
rect 54402 87502 54414 87554
rect 59154 87502 59166 87554
rect 59218 87502 59230 87554
rect 64306 87502 64318 87554
rect 64370 87502 64382 87554
rect 72258 87502 72270 87554
rect 72322 87502 72334 87554
rect 89506 87502 89518 87554
rect 89570 87502 89582 87554
rect 87278 87490 87330 87502
rect 1710 87442 1762 87454
rect 55582 87442 55634 87454
rect 54226 87390 54238 87442
rect 54290 87390 54302 87442
rect 1710 87378 1762 87390
rect 55582 87378 55634 87390
rect 56030 87442 56082 87454
rect 65326 87442 65378 87454
rect 70702 87442 70754 87454
rect 95118 87442 95170 87454
rect 59042 87390 59054 87442
rect 59106 87390 59118 87442
rect 59938 87390 59950 87442
rect 60002 87390 60014 87442
rect 64530 87390 64542 87442
rect 64594 87390 64606 87442
rect 67442 87390 67454 87442
rect 67506 87390 67518 87442
rect 72482 87390 72494 87442
rect 72546 87390 72558 87442
rect 87042 87390 87054 87442
rect 87106 87390 87118 87442
rect 94546 87390 94558 87442
rect 94610 87390 94622 87442
rect 56030 87378 56082 87390
rect 65326 87378 65378 87390
rect 70702 87378 70754 87390
rect 95118 87378 95170 87390
rect 55022 87330 55074 87342
rect 55022 87266 55074 87278
rect 57486 87330 57538 87342
rect 73278 87330 73330 87342
rect 60610 87278 60622 87330
rect 60674 87278 60686 87330
rect 62738 87278 62750 87330
rect 62802 87278 62814 87330
rect 68114 87278 68126 87330
rect 68178 87278 68190 87330
rect 70242 87278 70254 87330
rect 70306 87278 70318 87330
rect 57486 87266 57538 87278
rect 73278 87266 73330 87278
rect 73726 87330 73778 87342
rect 73726 87266 73778 87278
rect 74510 87330 74562 87342
rect 74510 87266 74562 87278
rect 75070 87330 75122 87342
rect 75070 87266 75122 87278
rect 75518 87330 75570 87342
rect 75518 87266 75570 87278
rect 53230 87218 53282 87230
rect 53230 87154 53282 87166
rect 53566 87218 53618 87230
rect 53566 87154 53618 87166
rect 58382 87218 58434 87230
rect 58382 87154 58434 87166
rect 63422 87218 63474 87230
rect 63422 87154 63474 87166
rect 63758 87218 63810 87230
rect 63758 87154 63810 87166
rect 71374 87218 71426 87230
rect 71374 87154 71426 87166
rect 71710 87218 71762 87230
rect 71710 87154 71762 87166
rect 1344 87050 98560 87084
rect 1344 86998 4478 87050
rect 4530 86998 4582 87050
rect 4634 86998 4686 87050
rect 4738 86998 35198 87050
rect 35250 86998 35302 87050
rect 35354 86998 35406 87050
rect 35458 86998 65918 87050
rect 65970 86998 66022 87050
rect 66074 86998 66126 87050
rect 66178 86998 96638 87050
rect 96690 86998 96742 87050
rect 96794 86998 96846 87050
rect 96898 86998 98560 87050
rect 1344 86964 98560 86998
rect 81790 86882 81842 86894
rect 81790 86818 81842 86830
rect 87614 86882 87666 86894
rect 87614 86818 87666 86830
rect 60622 86770 60674 86782
rect 57138 86718 57150 86770
rect 57202 86718 57214 86770
rect 59266 86718 59278 86770
rect 59330 86718 59342 86770
rect 60622 86706 60674 86718
rect 62190 86770 62242 86782
rect 73166 86770 73218 86782
rect 65762 86718 65774 86770
rect 65826 86718 65838 86770
rect 74722 86718 74734 86770
rect 74786 86718 74798 86770
rect 62190 86706 62242 86718
rect 73166 86706 73218 86718
rect 52558 86658 52610 86670
rect 52558 86594 52610 86606
rect 53902 86658 53954 86670
rect 69806 86658 69858 86670
rect 54674 86606 54686 86658
rect 54738 86606 54750 86658
rect 55570 86606 55582 86658
rect 55634 86606 55646 86658
rect 56466 86606 56478 86658
rect 56530 86606 56542 86658
rect 60050 86606 60062 86658
rect 60114 86606 60126 86658
rect 61618 86606 61630 86658
rect 61682 86606 61694 86658
rect 62962 86606 62974 86658
rect 63026 86606 63038 86658
rect 53902 86594 53954 86606
rect 69806 86594 69858 86606
rect 71710 86658 71762 86670
rect 71710 86594 71762 86606
rect 73726 86658 73778 86670
rect 87950 86658 88002 86670
rect 74386 86606 74398 86658
rect 74450 86606 74462 86658
rect 77858 86606 77870 86658
rect 77922 86606 77934 86658
rect 73726 86594 73778 86606
rect 87950 86594 88002 86606
rect 61406 86546 61458 86558
rect 68238 86546 68290 86558
rect 54450 86494 54462 86546
rect 54514 86494 54526 86546
rect 63634 86494 63646 86546
rect 63698 86494 63710 86546
rect 61406 86482 61458 86494
rect 68238 86482 68290 86494
rect 68574 86546 68626 86558
rect 71374 86546 71426 86558
rect 75742 86546 75794 86558
rect 70130 86494 70142 86546
rect 70194 86494 70206 86546
rect 70354 86494 70366 86546
rect 70418 86494 70430 86546
rect 71922 86494 71934 86546
rect 71986 86494 71998 86546
rect 72258 86494 72270 86546
rect 72322 86494 72334 86546
rect 68574 86482 68626 86494
rect 71374 86482 71426 86494
rect 75742 86482 75794 86494
rect 81902 86546 81954 86558
rect 81902 86482 81954 86494
rect 82462 86546 82514 86558
rect 82462 86482 82514 86494
rect 86494 86546 86546 86558
rect 91534 86546 91586 86558
rect 88162 86494 88174 86546
rect 88226 86494 88238 86546
rect 88722 86494 88734 86546
rect 88786 86494 88798 86546
rect 86494 86482 86546 86494
rect 91534 86482 91586 86494
rect 91870 86546 91922 86558
rect 91870 86482 91922 86494
rect 95566 86546 95618 86558
rect 95566 86482 95618 86494
rect 52222 86434 52274 86446
rect 52222 86370 52274 86382
rect 53566 86434 53618 86446
rect 53566 86370 53618 86382
rect 55358 86434 55410 86446
rect 55358 86370 55410 86382
rect 59838 86434 59890 86446
rect 59838 86370 59890 86382
rect 66334 86434 66386 86446
rect 66334 86370 66386 86382
rect 66670 86434 66722 86446
rect 66670 86370 66722 86382
rect 69470 86434 69522 86446
rect 69470 86370 69522 86382
rect 75406 86434 75458 86446
rect 75406 86370 75458 86382
rect 76526 86434 76578 86446
rect 76526 86370 76578 86382
rect 77310 86434 77362 86446
rect 77310 86370 77362 86382
rect 78094 86434 78146 86446
rect 78094 86370 78146 86382
rect 78654 86434 78706 86446
rect 78654 86370 78706 86382
rect 79662 86434 79714 86446
rect 79662 86370 79714 86382
rect 81230 86434 81282 86446
rect 81230 86370 81282 86382
rect 81790 86434 81842 86446
rect 81790 86370 81842 86382
rect 82574 86434 82626 86446
rect 82574 86370 82626 86382
rect 82798 86434 82850 86446
rect 82798 86370 82850 86382
rect 83134 86434 83186 86446
rect 83134 86370 83186 86382
rect 86158 86434 86210 86446
rect 86158 86370 86210 86382
rect 87054 86434 87106 86446
rect 87054 86370 87106 86382
rect 89294 86434 89346 86446
rect 89294 86370 89346 86382
rect 95902 86434 95954 86446
rect 95902 86370 95954 86382
rect 1344 86266 98560 86300
rect 1344 86214 19838 86266
rect 19890 86214 19942 86266
rect 19994 86214 20046 86266
rect 20098 86214 50558 86266
rect 50610 86214 50662 86266
rect 50714 86214 50766 86266
rect 50818 86214 81278 86266
rect 81330 86214 81382 86266
rect 81434 86214 81486 86266
rect 81538 86214 98560 86266
rect 1344 86180 98560 86214
rect 55470 86098 55522 86110
rect 55470 86034 55522 86046
rect 72718 86098 72770 86110
rect 72718 86034 72770 86046
rect 73390 86098 73442 86110
rect 73390 86034 73442 86046
rect 79214 86098 79266 86110
rect 79214 86034 79266 86046
rect 95902 85986 95954 85998
rect 56578 85934 56590 85986
rect 56642 85934 56654 85986
rect 58258 85934 58270 85986
rect 58322 85934 58334 85986
rect 75282 85934 75294 85986
rect 75346 85934 75358 85986
rect 78194 85934 78206 85986
rect 78258 85934 78270 85986
rect 78642 85934 78654 85986
rect 78706 85934 78718 85986
rect 87714 85934 87726 85986
rect 87778 85934 87790 85986
rect 95902 85922 95954 85934
rect 95566 85874 95618 85886
rect 51202 85822 51214 85874
rect 51266 85822 51278 85874
rect 56466 85822 56478 85874
rect 56530 85822 56542 85874
rect 57586 85822 57598 85874
rect 57650 85822 57662 85874
rect 63074 85822 63086 85874
rect 63138 85822 63150 85874
rect 63858 85822 63870 85874
rect 63922 85822 63934 85874
rect 66434 85822 66446 85874
rect 66498 85822 66510 85874
rect 74610 85822 74622 85874
rect 74674 85822 74686 85874
rect 84242 85822 84254 85874
rect 84306 85822 84318 85874
rect 88386 85822 88398 85874
rect 88450 85822 88462 85874
rect 93538 85822 93550 85874
rect 93602 85822 93614 85874
rect 95566 85810 95618 85822
rect 54574 85762 54626 85774
rect 51874 85710 51886 85762
rect 51938 85710 51950 85762
rect 54002 85710 54014 85762
rect 54066 85710 54078 85762
rect 54574 85698 54626 85710
rect 55806 85762 55858 85774
rect 64318 85762 64370 85774
rect 60386 85710 60398 85762
rect 60450 85710 60462 85762
rect 60946 85710 60958 85762
rect 61010 85710 61022 85762
rect 55806 85698 55858 85710
rect 64318 85698 64370 85710
rect 65438 85762 65490 85774
rect 71710 85762 71762 85774
rect 78878 85762 78930 85774
rect 69458 85710 69470 85762
rect 69522 85710 69534 85762
rect 73826 85710 73838 85762
rect 73890 85710 73902 85762
rect 77410 85710 77422 85762
rect 77474 85710 77486 85762
rect 65438 85698 65490 85710
rect 71710 85698 71762 85710
rect 78878 85698 78930 85710
rect 79774 85762 79826 85774
rect 79774 85698 79826 85710
rect 80446 85762 80498 85774
rect 84814 85762 84866 85774
rect 89182 85762 89234 85774
rect 81330 85710 81342 85762
rect 81394 85710 81406 85762
rect 83458 85710 83470 85762
rect 83522 85710 83534 85762
rect 85586 85710 85598 85762
rect 85650 85710 85662 85762
rect 90626 85710 90638 85762
rect 90690 85710 90702 85762
rect 92754 85710 92766 85762
rect 92818 85710 92830 85762
rect 80446 85698 80498 85710
rect 84814 85698 84866 85710
rect 89182 85698 89234 85710
rect 1344 85482 98560 85516
rect 1344 85430 4478 85482
rect 4530 85430 4582 85482
rect 4634 85430 4686 85482
rect 4738 85430 35198 85482
rect 35250 85430 35302 85482
rect 35354 85430 35406 85482
rect 35458 85430 65918 85482
rect 65970 85430 66022 85482
rect 66074 85430 66126 85482
rect 66178 85430 96638 85482
rect 96690 85430 96742 85482
rect 96794 85430 96846 85482
rect 96898 85430 98560 85482
rect 1344 85396 98560 85430
rect 59390 85314 59442 85326
rect 59390 85250 59442 85262
rect 59726 85314 59778 85326
rect 59726 85250 59778 85262
rect 74958 85314 75010 85326
rect 74958 85250 75010 85262
rect 75294 85314 75346 85326
rect 75294 85250 75346 85262
rect 88846 85314 88898 85326
rect 88846 85250 88898 85262
rect 91198 85314 91250 85326
rect 91198 85250 91250 85262
rect 57710 85202 57762 85214
rect 55122 85150 55134 85202
rect 55186 85150 55198 85202
rect 57250 85150 57262 85202
rect 57314 85150 57326 85202
rect 57710 85138 57762 85150
rect 60286 85202 60338 85214
rect 73166 85202 73218 85214
rect 89182 85202 89234 85214
rect 62626 85150 62638 85202
rect 62690 85150 62702 85202
rect 64754 85150 64766 85202
rect 64818 85150 64830 85202
rect 72258 85150 72270 85202
rect 72322 85150 72334 85202
rect 86034 85150 86046 85202
rect 86098 85150 86110 85202
rect 88162 85150 88174 85202
rect 88226 85150 88238 85202
rect 95666 85150 95678 85202
rect 95730 85150 95742 85202
rect 97794 85150 97806 85202
rect 97858 85150 97870 85202
rect 60286 85138 60338 85150
rect 73166 85138 73218 85150
rect 89182 85138 89234 85150
rect 52558 85090 52610 85102
rect 66558 85090 66610 85102
rect 68350 85090 68402 85102
rect 91534 85090 91586 85102
rect 54450 85038 54462 85090
rect 54514 85038 54526 85090
rect 61506 85038 61518 85090
rect 61570 85038 61582 85090
rect 65538 85038 65550 85090
rect 65602 85038 65614 85090
rect 67106 85038 67118 85090
rect 67170 85038 67182 85090
rect 69458 85038 69470 85090
rect 69522 85038 69534 85090
rect 74050 85038 74062 85090
rect 74114 85038 74126 85090
rect 82562 85038 82574 85090
rect 82626 85038 82638 85090
rect 85362 85038 85374 85090
rect 85426 85038 85438 85090
rect 89618 85038 89630 85090
rect 89682 85038 89694 85090
rect 92194 85038 92206 85090
rect 92258 85038 92270 85090
rect 93426 85038 93438 85090
rect 93490 85038 93502 85090
rect 94882 85038 94894 85090
rect 94946 85038 94958 85090
rect 52558 85026 52610 85038
rect 66558 85026 66610 85038
rect 68350 85026 68402 85038
rect 91534 85026 91586 85038
rect 52222 84978 52274 84990
rect 61742 84978 61794 84990
rect 93214 84978 93266 84990
rect 58706 84926 58718 84978
rect 58770 84926 58782 84978
rect 59042 84926 59054 84978
rect 59106 84926 59118 84978
rect 67218 84926 67230 84978
rect 67282 84926 67294 84978
rect 70130 84926 70142 84978
rect 70194 84926 70206 84978
rect 75618 84926 75630 84978
rect 75682 84926 75694 84978
rect 76066 84926 76078 84978
rect 76130 84926 76142 84978
rect 78754 84926 78766 84978
rect 78818 84926 78830 84978
rect 89730 84926 89742 84978
rect 89794 84926 89806 84978
rect 92306 84926 92318 84978
rect 92370 84926 92382 84978
rect 52222 84914 52274 84926
rect 61742 84914 61794 84926
rect 93214 84914 93266 84926
rect 53790 84866 53842 84878
rect 53790 84802 53842 84814
rect 66222 84866 66274 84878
rect 66222 84802 66274 84814
rect 68014 84866 68066 84878
rect 68014 84802 68066 84814
rect 72830 84866 72882 84878
rect 72830 84802 72882 84814
rect 74286 84866 74338 84878
rect 74286 84802 74338 84814
rect 83022 84866 83074 84878
rect 83022 84802 83074 84814
rect 83470 84866 83522 84878
rect 83470 84802 83522 84814
rect 90526 84866 90578 84878
rect 90526 84802 90578 84814
rect 94446 84866 94498 84878
rect 94446 84802 94498 84814
rect 1344 84698 98560 84732
rect 1344 84646 19838 84698
rect 19890 84646 19942 84698
rect 19994 84646 20046 84698
rect 20098 84646 50558 84698
rect 50610 84646 50662 84698
rect 50714 84646 50766 84698
rect 50818 84646 81278 84698
rect 81330 84646 81382 84698
rect 81434 84646 81486 84698
rect 81538 84646 98560 84698
rect 1344 84612 98560 84646
rect 65774 84530 65826 84542
rect 65774 84466 65826 84478
rect 90526 84530 90578 84542
rect 90526 84466 90578 84478
rect 95230 84530 95282 84542
rect 95230 84466 95282 84478
rect 84926 84418 84978 84430
rect 89294 84418 89346 84430
rect 51762 84366 51774 84418
rect 51826 84366 51838 84418
rect 60610 84366 60622 84418
rect 60674 84366 60686 84418
rect 67106 84366 67118 84418
rect 67170 84366 67182 84418
rect 71026 84366 71038 84418
rect 71090 84366 71102 84418
rect 74274 84366 74286 84418
rect 74338 84366 74350 84418
rect 78082 84366 78094 84418
rect 78146 84366 78158 84418
rect 87714 84366 87726 84418
rect 87778 84366 87790 84418
rect 95778 84366 95790 84418
rect 95842 84366 95854 84418
rect 96338 84366 96350 84418
rect 96402 84366 96414 84418
rect 84926 84354 84978 84366
rect 89294 84354 89346 84366
rect 64318 84306 64370 84318
rect 71934 84306 71986 84318
rect 51090 84254 51102 84306
rect 51154 84254 51166 84306
rect 58818 84254 58830 84306
rect 58882 84254 58894 84306
rect 66322 84254 66334 84306
rect 66386 84254 66398 84306
rect 71250 84254 71262 84306
rect 71314 84254 71326 84306
rect 64318 84242 64370 84254
rect 71934 84242 71986 84254
rect 72494 84306 72546 84318
rect 85038 84306 85090 84318
rect 90190 84306 90242 84318
rect 95566 84306 95618 84318
rect 73602 84254 73614 84306
rect 73666 84254 73678 84306
rect 77410 84254 77422 84306
rect 77474 84254 77486 84306
rect 81442 84254 81454 84306
rect 81506 84254 81518 84306
rect 88498 84254 88510 84306
rect 88562 84254 88574 84306
rect 89506 84254 89518 84306
rect 89570 84254 89582 84306
rect 94434 84254 94446 84306
rect 94498 84254 94510 84306
rect 72494 84242 72546 84254
rect 85038 84242 85090 84254
rect 90190 84242 90242 84254
rect 95566 84242 95618 84254
rect 54462 84194 54514 84206
rect 53890 84142 53902 84194
rect 53954 84142 53966 84194
rect 54462 84130 54514 84142
rect 54798 84194 54850 84206
rect 54798 84130 54850 84142
rect 57374 84194 57426 84206
rect 90974 84194 91026 84206
rect 69234 84142 69246 84194
rect 69298 84142 69310 84194
rect 76402 84142 76414 84194
rect 76466 84142 76478 84194
rect 80210 84142 80222 84194
rect 80274 84142 80286 84194
rect 82114 84142 82126 84194
rect 82178 84142 82190 84194
rect 84242 84142 84254 84194
rect 84306 84142 84318 84194
rect 85586 84142 85598 84194
rect 85650 84142 85662 84194
rect 91522 84142 91534 84194
rect 91586 84142 91598 84194
rect 93650 84142 93662 84194
rect 93714 84142 93726 84194
rect 57374 84130 57426 84142
rect 90974 84130 91026 84142
rect 70142 84082 70194 84094
rect 70142 84018 70194 84030
rect 70478 84082 70530 84094
rect 70478 84018 70530 84030
rect 84926 84082 84978 84094
rect 84926 84018 84978 84030
rect 1344 83914 98560 83948
rect 1344 83862 4478 83914
rect 4530 83862 4582 83914
rect 4634 83862 4686 83914
rect 4738 83862 35198 83914
rect 35250 83862 35302 83914
rect 35354 83862 35406 83914
rect 35458 83862 65918 83914
rect 65970 83862 66022 83914
rect 66074 83862 66126 83914
rect 66178 83862 96638 83914
rect 96690 83862 96742 83914
rect 96794 83862 96846 83914
rect 96898 83862 98560 83914
rect 1344 83828 98560 83862
rect 63422 83746 63474 83758
rect 63422 83682 63474 83694
rect 74286 83746 74338 83758
rect 74286 83682 74338 83694
rect 74622 83746 74674 83758
rect 74622 83682 74674 83694
rect 83694 83746 83746 83758
rect 83694 83682 83746 83694
rect 88286 83746 88338 83758
rect 88286 83682 88338 83694
rect 88622 83746 88674 83758
rect 88622 83682 88674 83694
rect 91198 83746 91250 83758
rect 91198 83682 91250 83694
rect 65102 83634 65154 83646
rect 65102 83570 65154 83582
rect 67678 83634 67730 83646
rect 67678 83570 67730 83582
rect 79550 83634 79602 83646
rect 90526 83634 90578 83646
rect 83010 83582 83022 83634
rect 83074 83582 83086 83634
rect 79550 83570 79602 83582
rect 90526 83570 90578 83582
rect 94334 83634 94386 83646
rect 95666 83582 95678 83634
rect 95730 83582 95742 83634
rect 97794 83582 97806 83634
rect 97858 83582 97870 83634
rect 94334 83570 94386 83582
rect 53678 83522 53730 83534
rect 63758 83522 63810 83534
rect 69694 83522 69746 83534
rect 57922 83470 57934 83522
rect 57986 83470 57998 83522
rect 64418 83470 64430 83522
rect 64482 83470 64494 83522
rect 53678 83458 53730 83470
rect 63758 83458 63810 83470
rect 69694 83458 69746 83470
rect 70590 83522 70642 83534
rect 73166 83522 73218 83534
rect 78206 83522 78258 83534
rect 91534 83522 91586 83534
rect 72706 83470 72718 83522
rect 72770 83470 72782 83522
rect 77522 83470 77534 83522
rect 77586 83470 77598 83522
rect 80210 83470 80222 83522
rect 80274 83470 80286 83522
rect 92194 83470 92206 83522
rect 92258 83470 92270 83522
rect 93314 83470 93326 83522
rect 93378 83470 93390 83522
rect 94882 83470 94894 83522
rect 94946 83470 94958 83522
rect 70590 83458 70642 83470
rect 73166 83458 73218 83470
rect 78206 83458 78258 83470
rect 91534 83458 91586 83470
rect 54462 83410 54514 83422
rect 69358 83410 69410 83422
rect 64530 83358 64542 83410
rect 64594 83358 64606 83410
rect 54462 83346 54514 83358
rect 69358 83346 69410 83358
rect 70254 83410 70306 83422
rect 76414 83410 76466 83422
rect 78542 83410 78594 83422
rect 83582 83410 83634 83422
rect 93550 83410 93602 83422
rect 74946 83358 74958 83410
rect 75010 83358 75022 83410
rect 75394 83358 75406 83410
rect 75458 83358 75470 83410
rect 77410 83358 77422 83410
rect 77474 83358 77486 83410
rect 80882 83358 80894 83410
rect 80946 83358 80958 83410
rect 88834 83358 88846 83410
rect 88898 83358 88910 83410
rect 89394 83358 89406 83410
rect 89458 83358 89470 83410
rect 92306 83358 92318 83410
rect 92370 83358 92382 83410
rect 70254 83346 70306 83358
rect 76414 83346 76466 83358
rect 78542 83346 78594 83358
rect 83582 83346 83634 83358
rect 93550 83346 93602 83358
rect 52670 83298 52722 83310
rect 52670 83234 52722 83246
rect 53342 83298 53394 83310
rect 53342 83234 53394 83246
rect 53566 83298 53618 83310
rect 53566 83234 53618 83246
rect 54126 83298 54178 83310
rect 54126 83234 54178 83246
rect 54350 83298 54402 83310
rect 54350 83234 54402 83246
rect 54910 83298 54962 83310
rect 54910 83234 54962 83246
rect 56926 83298 56978 83310
rect 56926 83234 56978 83246
rect 58158 83298 58210 83310
rect 58158 83234 58210 83246
rect 71598 83298 71650 83310
rect 71598 83234 71650 83246
rect 73614 83298 73666 83310
rect 73614 83234 73666 83246
rect 76078 83298 76130 83310
rect 76078 83234 76130 83246
rect 79214 83298 79266 83310
rect 79214 83234 79266 83246
rect 83694 83298 83746 83310
rect 83694 83234 83746 83246
rect 84366 83298 84418 83310
rect 84366 83234 84418 83246
rect 85262 83298 85314 83310
rect 85262 83234 85314 83246
rect 85710 83298 85762 83310
rect 85710 83234 85762 83246
rect 87614 83298 87666 83310
rect 87614 83234 87666 83246
rect 1344 83130 98560 83164
rect 1344 83078 19838 83130
rect 19890 83078 19942 83130
rect 19994 83078 20046 83130
rect 20098 83078 50558 83130
rect 50610 83078 50662 83130
rect 50714 83078 50766 83130
rect 50818 83078 81278 83130
rect 81330 83078 81382 83130
rect 81434 83078 81486 83130
rect 81538 83078 98560 83130
rect 1344 83044 98560 83078
rect 60846 82962 60898 82974
rect 60846 82898 60898 82910
rect 63422 82962 63474 82974
rect 63422 82898 63474 82910
rect 74846 82962 74898 82974
rect 74846 82898 74898 82910
rect 78766 82962 78818 82974
rect 78766 82898 78818 82910
rect 80446 82962 80498 82974
rect 80446 82898 80498 82910
rect 61630 82850 61682 82862
rect 58258 82798 58270 82850
rect 58322 82798 58334 82850
rect 61630 82786 61682 82798
rect 63758 82850 63810 82862
rect 76178 82798 76190 82850
rect 76242 82798 76254 82850
rect 82674 82798 82686 82850
rect 82738 82798 82750 82850
rect 63758 82786 63810 82798
rect 61966 82738 62018 82750
rect 80334 82738 80386 82750
rect 52882 82686 52894 82738
rect 52946 82686 52958 82738
rect 57586 82686 57598 82738
rect 57650 82686 57662 82738
rect 75506 82686 75518 82738
rect 75570 82686 75582 82738
rect 82002 82686 82014 82738
rect 82066 82686 82078 82738
rect 92642 82686 92654 82738
rect 92706 82686 92718 82738
rect 61966 82674 62018 82686
rect 80334 82674 80386 82686
rect 69470 82626 69522 82638
rect 54114 82574 54126 82626
rect 54178 82574 54190 82626
rect 60386 82574 60398 82626
rect 60450 82574 60462 82626
rect 69470 82562 69522 82574
rect 69918 82626 69970 82638
rect 69918 82562 69970 82574
rect 73838 82626 73890 82638
rect 81454 82626 81506 82638
rect 85262 82626 85314 82638
rect 78306 82574 78318 82626
rect 78370 82574 78382 82626
rect 84802 82574 84814 82626
rect 84866 82574 84878 82626
rect 73838 82562 73890 82574
rect 81454 82562 81506 82574
rect 85262 82562 85314 82574
rect 85822 82626 85874 82638
rect 85822 82562 85874 82574
rect 86158 82626 86210 82638
rect 86158 82562 86210 82574
rect 86606 82626 86658 82638
rect 86606 82562 86658 82574
rect 90638 82626 90690 82638
rect 94882 82574 94894 82626
rect 94946 82574 94958 82626
rect 90638 82562 90690 82574
rect 80446 82514 80498 82526
rect 85698 82462 85710 82514
rect 85762 82511 85774 82514
rect 86706 82511 86718 82514
rect 85762 82465 86718 82511
rect 85762 82462 85774 82465
rect 86706 82462 86718 82465
rect 86770 82462 86782 82514
rect 80446 82450 80498 82462
rect 1344 82346 98560 82380
rect 1344 82294 4478 82346
rect 4530 82294 4582 82346
rect 4634 82294 4686 82346
rect 4738 82294 35198 82346
rect 35250 82294 35302 82346
rect 35354 82294 35406 82346
rect 35458 82294 65918 82346
rect 65970 82294 66022 82346
rect 66074 82294 66126 82346
rect 66178 82294 96638 82346
rect 96690 82294 96742 82346
rect 96794 82294 96846 82346
rect 96898 82294 98560 82346
rect 1344 82260 98560 82294
rect 58606 82178 58658 82190
rect 58606 82114 58658 82126
rect 62302 82178 62354 82190
rect 62302 82114 62354 82126
rect 93326 82178 93378 82190
rect 93326 82114 93378 82126
rect 95230 82178 95282 82190
rect 95230 82114 95282 82126
rect 63982 82066 64034 82078
rect 75406 82066 75458 82078
rect 52658 82014 52670 82066
rect 52722 82014 52734 82066
rect 57026 82014 57038 82066
rect 57090 82014 57102 82066
rect 73266 82014 73278 82066
rect 73330 82014 73342 82066
rect 63982 82002 64034 82014
rect 75406 82002 75458 82014
rect 77870 82066 77922 82078
rect 77870 82002 77922 82014
rect 97358 82066 97410 82078
rect 97358 82002 97410 82014
rect 58942 81954 58994 81966
rect 62638 81954 62690 81966
rect 81118 81954 81170 81966
rect 49746 81902 49758 81954
rect 49810 81902 49822 81954
rect 54114 81902 54126 81954
rect 54178 81902 54190 81954
rect 59714 81902 59726 81954
rect 59778 81902 59790 81954
rect 63410 81902 63422 81954
rect 63474 81902 63486 81954
rect 58942 81890 58994 81902
rect 62638 81890 62690 81902
rect 81118 81890 81170 81902
rect 81454 81954 81506 81966
rect 81454 81890 81506 81902
rect 82686 81954 82738 81966
rect 82686 81890 82738 81902
rect 83022 81954 83074 81966
rect 83022 81890 83074 81902
rect 83918 81954 83970 81966
rect 93662 81954 93714 81966
rect 86706 81902 86718 81954
rect 86770 81902 86782 81954
rect 83918 81890 83970 81902
rect 93662 81890 93714 81902
rect 95566 81954 95618 81966
rect 96226 81902 96238 81954
rect 96290 81902 96302 81954
rect 95566 81890 95618 81902
rect 68014 81842 68066 81854
rect 50530 81790 50542 81842
rect 50594 81790 50606 81842
rect 54898 81790 54910 81842
rect 54962 81790 54974 81842
rect 59490 81790 59502 81842
rect 59554 81790 59566 81842
rect 63186 81790 63198 81842
rect 63250 81790 63262 81842
rect 68014 81778 68066 81790
rect 72830 81842 72882 81854
rect 72830 81778 72882 81790
rect 83582 81842 83634 81854
rect 87602 81790 87614 81842
rect 87666 81790 87678 81842
rect 93874 81790 93886 81842
rect 93938 81790 93950 81842
rect 94210 81790 94222 81842
rect 94274 81790 94286 81842
rect 96338 81790 96350 81842
rect 96402 81790 96414 81842
rect 83582 81778 83634 81790
rect 53342 81730 53394 81742
rect 53342 81666 53394 81678
rect 60286 81730 60338 81742
rect 60286 81666 60338 81678
rect 64430 81730 64482 81742
rect 64430 81666 64482 81678
rect 68126 81730 68178 81742
rect 68126 81666 68178 81678
rect 68350 81730 68402 81742
rect 68350 81666 68402 81678
rect 69806 81730 69858 81742
rect 69806 81666 69858 81678
rect 70366 81730 70418 81742
rect 70366 81666 70418 81678
rect 73838 81730 73890 81742
rect 73838 81666 73890 81678
rect 74286 81730 74338 81742
rect 74286 81666 74338 81678
rect 74846 81730 74898 81742
rect 74846 81666 74898 81678
rect 76526 81730 76578 81742
rect 76526 81666 76578 81678
rect 77310 81730 77362 81742
rect 77310 81666 77362 81678
rect 80670 81730 80722 81742
rect 80670 81666 80722 81678
rect 81342 81730 81394 81742
rect 81342 81666 81394 81678
rect 82014 81730 82066 81742
rect 82014 81666 82066 81678
rect 82910 81730 82962 81742
rect 82910 81666 82962 81678
rect 83694 81730 83746 81742
rect 83694 81666 83746 81678
rect 84366 81730 84418 81742
rect 84366 81666 84418 81678
rect 90974 81730 91026 81742
rect 90974 81666 91026 81678
rect 92430 81730 92482 81742
rect 92430 81666 92482 81678
rect 96910 81730 96962 81742
rect 96910 81666 96962 81678
rect 97806 81730 97858 81742
rect 97806 81666 97858 81678
rect 1344 81562 98560 81596
rect 1344 81510 19838 81562
rect 19890 81510 19942 81562
rect 19994 81510 20046 81562
rect 20098 81510 50558 81562
rect 50610 81510 50662 81562
rect 50714 81510 50766 81562
rect 50818 81510 81278 81562
rect 81330 81510 81382 81562
rect 81434 81510 81486 81562
rect 81538 81510 98560 81562
rect 1344 81476 98560 81510
rect 50766 81394 50818 81406
rect 50766 81330 50818 81342
rect 56590 81394 56642 81406
rect 56590 81330 56642 81342
rect 69694 81394 69746 81406
rect 69694 81330 69746 81342
rect 73838 81394 73890 81406
rect 73838 81330 73890 81342
rect 74510 81394 74562 81406
rect 74510 81330 74562 81342
rect 75070 81394 75122 81406
rect 75070 81330 75122 81342
rect 80558 81394 80610 81406
rect 80558 81330 80610 81342
rect 92206 81394 92258 81406
rect 92206 81330 92258 81342
rect 50206 81282 50258 81294
rect 50206 81218 50258 81230
rect 50318 81282 50370 81294
rect 50318 81218 50370 81230
rect 50990 81282 51042 81294
rect 55246 81282 55298 81294
rect 52434 81230 52446 81282
rect 52498 81230 52510 81282
rect 50990 81218 51042 81230
rect 55246 81218 55298 81230
rect 56030 81282 56082 81294
rect 63982 81282 64034 81294
rect 81454 81282 81506 81294
rect 61282 81230 61294 81282
rect 61346 81230 61358 81282
rect 68450 81230 68462 81282
rect 68514 81230 68526 81282
rect 56030 81218 56082 81230
rect 63982 81218 64034 81230
rect 81454 81218 81506 81230
rect 82350 81282 82402 81294
rect 82350 81218 82402 81230
rect 83134 81282 83186 81294
rect 83134 81218 83186 81230
rect 83246 81282 83298 81294
rect 83246 81218 83298 81230
rect 85262 81282 85314 81294
rect 86258 81230 86270 81282
rect 86322 81230 86334 81282
rect 93538 81230 93550 81282
rect 93602 81230 93614 81282
rect 93762 81230 93774 81282
rect 93826 81230 93838 81282
rect 95778 81230 95790 81282
rect 95842 81230 95854 81282
rect 96114 81230 96126 81282
rect 96178 81230 96190 81282
rect 85262 81218 85314 81230
rect 51102 81170 51154 81182
rect 55022 81170 55074 81182
rect 51650 81118 51662 81170
rect 51714 81118 51726 81170
rect 51102 81106 51154 81118
rect 55022 81106 55074 81118
rect 55358 81170 55410 81182
rect 55358 81106 55410 81118
rect 55806 81170 55858 81182
rect 55806 81106 55858 81118
rect 56142 81170 56194 81182
rect 71486 81170 71538 81182
rect 60610 81118 60622 81170
rect 60674 81118 60686 81170
rect 64194 81118 64206 81170
rect 64258 81118 64270 81170
rect 69234 81118 69246 81170
rect 69298 81118 69310 81170
rect 56142 81106 56194 81118
rect 71486 81106 71538 81118
rect 72606 81170 72658 81182
rect 72606 81106 72658 81118
rect 73502 81170 73554 81182
rect 73502 81106 73554 81118
rect 74286 81170 74338 81182
rect 74286 81106 74338 81118
rect 74622 81170 74674 81182
rect 74622 81106 74674 81118
rect 80110 81170 80162 81182
rect 80110 81106 80162 81118
rect 81566 81170 81618 81182
rect 81566 81106 81618 81118
rect 82126 81170 82178 81182
rect 82126 81106 82178 81118
rect 82462 81170 82514 81182
rect 82462 81106 82514 81118
rect 82910 81170 82962 81182
rect 85698 81118 85710 81170
rect 85762 81118 85774 81170
rect 86034 81118 86046 81170
rect 86098 81118 86110 81170
rect 86818 81118 86830 81170
rect 86882 81118 86894 81170
rect 87490 81118 87502 81170
rect 87554 81118 87566 81170
rect 88386 81118 88398 81170
rect 88450 81118 88462 81170
rect 82910 81106 82962 81118
rect 57374 81058 57426 81070
rect 70142 81058 70194 81070
rect 54562 81006 54574 81058
rect 54626 81006 54638 81058
rect 63410 81006 63422 81058
rect 63474 81006 63486 81058
rect 66322 81006 66334 81058
rect 66386 81006 66398 81058
rect 57374 80994 57426 81006
rect 70142 80994 70194 81006
rect 70590 81058 70642 81070
rect 70590 80994 70642 81006
rect 71150 81058 71202 81070
rect 71150 80994 71202 81006
rect 72046 81058 72098 81070
rect 72046 80994 72098 81006
rect 83694 81058 83746 81070
rect 83694 80994 83746 81006
rect 84142 81058 84194 81070
rect 84142 80994 84194 81006
rect 84590 81058 84642 81070
rect 84590 80994 84642 81006
rect 93214 81058 93266 81070
rect 93214 80994 93266 81006
rect 94670 81058 94722 81070
rect 94670 80994 94722 81006
rect 95566 81058 95618 81070
rect 95566 80994 95618 81006
rect 97246 81058 97298 81070
rect 97246 80994 97298 81006
rect 50206 80946 50258 80958
rect 81454 80946 81506 80958
rect 71138 80894 71150 80946
rect 71202 80943 71214 80946
rect 71586 80943 71598 80946
rect 71202 80897 71598 80943
rect 71202 80894 71214 80897
rect 71586 80894 71598 80897
rect 71650 80943 71662 80946
rect 72034 80943 72046 80946
rect 71650 80897 72046 80943
rect 71650 80894 71662 80897
rect 72034 80894 72046 80897
rect 72098 80894 72110 80946
rect 50206 80882 50258 80894
rect 81454 80882 81506 80894
rect 92878 80946 92930 80958
rect 92878 80882 92930 80894
rect 95230 80946 95282 80958
rect 95230 80882 95282 80894
rect 1344 80778 98560 80812
rect 1344 80726 4478 80778
rect 4530 80726 4582 80778
rect 4634 80726 4686 80778
rect 4738 80726 35198 80778
rect 35250 80726 35302 80778
rect 35354 80726 35406 80778
rect 35458 80726 65918 80778
rect 65970 80726 66022 80778
rect 66074 80726 66126 80778
rect 66178 80726 96638 80778
rect 96690 80726 96742 80778
rect 96794 80726 96846 80778
rect 96898 80726 98560 80778
rect 1344 80692 98560 80726
rect 83582 80610 83634 80622
rect 85698 80558 85710 80610
rect 85762 80607 85774 80610
rect 86482 80607 86494 80610
rect 85762 80561 86494 80607
rect 85762 80558 85774 80561
rect 86482 80558 86494 80561
rect 86546 80558 86558 80610
rect 83582 80546 83634 80558
rect 85598 80498 85650 80510
rect 52322 80446 52334 80498
rect 52386 80446 52398 80498
rect 54226 80446 54238 80498
rect 54290 80446 54302 80498
rect 56354 80446 56366 80498
rect 56418 80446 56430 80498
rect 61394 80446 61406 80498
rect 61458 80446 61470 80498
rect 63522 80446 63534 80498
rect 63586 80446 63598 80498
rect 68562 80446 68574 80498
rect 68626 80446 68638 80498
rect 74498 80446 74510 80498
rect 74562 80446 74574 80498
rect 79538 80446 79550 80498
rect 79602 80446 79614 80498
rect 81666 80446 81678 80498
rect 81730 80446 81742 80498
rect 85598 80434 85650 80446
rect 86046 80498 86098 80510
rect 86046 80434 86098 80446
rect 86494 80498 86546 80510
rect 93102 80498 93154 80510
rect 88498 80446 88510 80498
rect 88562 80446 88574 80498
rect 86494 80434 86546 80446
rect 93102 80434 93154 80446
rect 93550 80498 93602 80510
rect 97794 80446 97806 80498
rect 97858 80446 97870 80498
rect 93550 80434 93602 80446
rect 56814 80386 56866 80398
rect 49522 80334 49534 80386
rect 49586 80334 49598 80386
rect 53442 80334 53454 80386
rect 53506 80334 53518 80386
rect 56814 80322 56866 80334
rect 57150 80386 57202 80398
rect 57150 80322 57202 80334
rect 57598 80386 57650 80398
rect 70030 80386 70082 80398
rect 64306 80334 64318 80386
rect 64370 80334 64382 80386
rect 65762 80334 65774 80386
rect 65826 80334 65838 80386
rect 57598 80322 57650 80334
rect 70030 80322 70082 80334
rect 70366 80386 70418 80398
rect 75294 80386 75346 80398
rect 82910 80386 82962 80398
rect 71698 80334 71710 80386
rect 71762 80334 71774 80386
rect 78866 80334 78878 80386
rect 78930 80334 78942 80386
rect 70366 80322 70418 80334
rect 75294 80322 75346 80334
rect 82910 80322 82962 80334
rect 84254 80386 84306 80398
rect 92418 80334 92430 80386
rect 92482 80334 92494 80386
rect 94882 80334 94894 80386
rect 94946 80334 94958 80386
rect 84254 80322 84306 80334
rect 57038 80274 57090 80286
rect 69470 80274 69522 80286
rect 50194 80222 50206 80274
rect 50258 80222 50270 80274
rect 66434 80222 66446 80274
rect 66498 80222 66510 80274
rect 57038 80210 57090 80222
rect 69470 80210 69522 80222
rect 69582 80274 69634 80286
rect 69582 80210 69634 80222
rect 70814 80274 70866 80286
rect 74958 80274 75010 80286
rect 72370 80222 72382 80274
rect 72434 80222 72446 80274
rect 70814 80210 70866 80222
rect 74958 80210 75010 80222
rect 75182 80274 75234 80286
rect 75182 80210 75234 80222
rect 83582 80274 83634 80286
rect 83582 80210 83634 80222
rect 83694 80274 83746 80286
rect 83694 80210 83746 80222
rect 94334 80274 94386 80286
rect 95666 80222 95678 80274
rect 95730 80222 95742 80274
rect 94334 80210 94386 80222
rect 64766 80162 64818 80174
rect 64766 80098 64818 80110
rect 69246 80162 69298 80174
rect 69246 80098 69298 80110
rect 70254 80162 70306 80174
rect 70254 80098 70306 80110
rect 75742 80162 75794 80174
rect 75742 80098 75794 80110
rect 76190 80162 76242 80174
rect 76190 80098 76242 80110
rect 82238 80162 82290 80174
rect 82238 80098 82290 80110
rect 82574 80162 82626 80174
rect 82574 80098 82626 80110
rect 82798 80162 82850 80174
rect 82798 80098 82850 80110
rect 84366 80162 84418 80174
rect 84366 80098 84418 80110
rect 84590 80162 84642 80174
rect 84590 80098 84642 80110
rect 85150 80162 85202 80174
rect 85150 80098 85202 80110
rect 1344 79994 98560 80028
rect 1344 79942 19838 79994
rect 19890 79942 19942 79994
rect 19994 79942 20046 79994
rect 20098 79942 50558 79994
rect 50610 79942 50662 79994
rect 50714 79942 50766 79994
rect 50818 79942 81278 79994
rect 81330 79942 81382 79994
rect 81434 79942 81486 79994
rect 81538 79942 98560 79994
rect 1344 79908 98560 79942
rect 52894 79826 52946 79838
rect 52894 79762 52946 79774
rect 53118 79826 53170 79838
rect 53118 79762 53170 79774
rect 53678 79826 53730 79838
rect 53678 79762 53730 79774
rect 54350 79826 54402 79838
rect 54350 79762 54402 79774
rect 55134 79826 55186 79838
rect 55134 79762 55186 79774
rect 55918 79826 55970 79838
rect 55918 79762 55970 79774
rect 56702 79826 56754 79838
rect 56702 79762 56754 79774
rect 63646 79826 63698 79838
rect 63646 79762 63698 79774
rect 64318 79826 64370 79838
rect 64318 79762 64370 79774
rect 70814 79826 70866 79838
rect 70814 79762 70866 79774
rect 71374 79826 71426 79838
rect 71374 79762 71426 79774
rect 72270 79826 72322 79838
rect 72270 79762 72322 79774
rect 80446 79826 80498 79838
rect 80446 79762 80498 79774
rect 84702 79826 84754 79838
rect 84702 79762 84754 79774
rect 89182 79826 89234 79838
rect 89182 79762 89234 79774
rect 89630 79826 89682 79838
rect 89630 79762 89682 79774
rect 97246 79826 97298 79838
rect 97246 79762 97298 79774
rect 53230 79714 53282 79726
rect 50306 79662 50318 79714
rect 50370 79662 50382 79714
rect 53230 79650 53282 79662
rect 54574 79714 54626 79726
rect 54574 79650 54626 79662
rect 55358 79714 55410 79726
rect 55358 79650 55410 79662
rect 55470 79714 55522 79726
rect 55470 79650 55522 79662
rect 57486 79714 57538 79726
rect 66446 79714 66498 79726
rect 80334 79714 80386 79726
rect 58482 79662 58494 79714
rect 58546 79662 58558 79714
rect 62738 79662 62750 79714
rect 62802 79662 62814 79714
rect 63074 79662 63086 79714
rect 63138 79662 63150 79714
rect 67442 79662 67454 79714
rect 67506 79662 67518 79714
rect 74162 79662 74174 79714
rect 74226 79662 74238 79714
rect 57486 79650 57538 79662
rect 66446 79650 66498 79662
rect 80334 79650 80386 79662
rect 80670 79714 80722 79726
rect 85262 79714 85314 79726
rect 95790 79714 95842 79726
rect 82114 79662 82126 79714
rect 82178 79662 82190 79714
rect 86258 79662 86270 79714
rect 86322 79662 86334 79714
rect 94546 79662 94558 79714
rect 94610 79662 94622 79714
rect 94882 79662 94894 79714
rect 94946 79662 94958 79714
rect 80670 79650 80722 79662
rect 85262 79650 85314 79662
rect 95790 79650 95842 79662
rect 96126 79714 96178 79726
rect 96126 79650 96178 79662
rect 54686 79602 54738 79614
rect 63310 79602 63362 79614
rect 68126 79602 68178 79614
rect 70478 79602 70530 79614
rect 97582 79602 97634 79614
rect 49522 79550 49534 79602
rect 49586 79550 49598 79602
rect 57922 79550 57934 79602
rect 57986 79550 57998 79602
rect 58258 79550 58270 79602
rect 58322 79550 58334 79602
rect 59042 79550 59054 79602
rect 59106 79550 59118 79602
rect 59490 79550 59502 79602
rect 59554 79550 59566 79602
rect 60498 79550 60510 79602
rect 60562 79550 60574 79602
rect 66770 79550 66782 79602
rect 66834 79550 66846 79602
rect 67218 79550 67230 79602
rect 67282 79550 67294 79602
rect 68674 79550 68686 79602
rect 68738 79550 68750 79602
rect 69570 79550 69582 79602
rect 69634 79550 69646 79602
rect 71586 79550 71598 79602
rect 71650 79550 71662 79602
rect 72482 79550 72494 79602
rect 72546 79550 72558 79602
rect 73490 79550 73502 79602
rect 73554 79550 73566 79602
rect 81442 79550 81454 79602
rect 81506 79550 81518 79602
rect 85586 79550 85598 79602
rect 85650 79550 85662 79602
rect 86034 79550 86046 79602
rect 86098 79550 86110 79602
rect 86818 79550 86830 79602
rect 86882 79550 86894 79602
rect 87490 79550 87502 79602
rect 87554 79550 87566 79602
rect 88386 79550 88398 79602
rect 88450 79550 88462 79602
rect 93314 79550 93326 79602
rect 93378 79550 93390 79602
rect 54686 79538 54738 79550
rect 63310 79538 63362 79550
rect 68126 79538 68178 79550
rect 70478 79538 70530 79550
rect 97582 79538 97634 79550
rect 61182 79490 61234 79502
rect 52434 79438 52446 79490
rect 52498 79438 52510 79490
rect 61182 79426 61234 79438
rect 61630 79490 61682 79502
rect 76750 79490 76802 79502
rect 76290 79438 76302 79490
rect 76354 79438 76366 79490
rect 61630 79426 61682 79438
rect 76750 79426 76802 79438
rect 77198 79490 77250 79502
rect 84242 79438 84254 79490
rect 84306 79438 84318 79490
rect 90402 79438 90414 79490
rect 90466 79438 90478 79490
rect 92530 79438 92542 79490
rect 92594 79438 92606 79490
rect 77198 79426 77250 79438
rect 93998 79378 94050 79390
rect 84466 79326 84478 79378
rect 84530 79375 84542 79378
rect 85026 79375 85038 79378
rect 84530 79329 85038 79375
rect 84530 79326 84542 79329
rect 85026 79326 85038 79329
rect 85090 79326 85102 79378
rect 93998 79314 94050 79326
rect 94334 79378 94386 79390
rect 94334 79314 94386 79326
rect 1344 79210 98560 79244
rect 1344 79158 4478 79210
rect 4530 79158 4582 79210
rect 4634 79158 4686 79210
rect 4738 79158 35198 79210
rect 35250 79158 35302 79210
rect 35354 79158 35406 79210
rect 35458 79158 65918 79210
rect 65970 79158 66022 79210
rect 66074 79158 66126 79210
rect 66178 79158 96638 79210
rect 96690 79158 96742 79210
rect 96794 79158 96846 79210
rect 96898 79158 98560 79210
rect 1344 79124 98560 79158
rect 54574 78930 54626 78942
rect 54574 78866 54626 78878
rect 57374 78930 57426 78942
rect 85262 78930 85314 78942
rect 67218 78878 67230 78930
rect 67282 78878 67294 78930
rect 73826 78878 73838 78930
rect 73890 78878 73902 78930
rect 80434 78878 80446 78930
rect 80498 78878 80510 78930
rect 57374 78866 57426 78878
rect 85262 78866 85314 78878
rect 88958 78930 89010 78942
rect 95666 78878 95678 78930
rect 95730 78878 95742 78930
rect 97794 78878 97806 78930
rect 97858 78878 97870 78930
rect 88958 78866 89010 78878
rect 52110 78818 52162 78830
rect 52110 78754 52162 78766
rect 52446 78818 52498 78830
rect 52446 78754 52498 78766
rect 53342 78818 53394 78830
rect 62302 78818 62354 78830
rect 68574 78818 68626 78830
rect 75966 78818 76018 78830
rect 83022 78818 83074 78830
rect 57810 78766 57822 78818
rect 57874 78766 57886 78818
rect 58258 78766 58270 78818
rect 58322 78766 58334 78818
rect 59378 78766 59390 78818
rect 59442 78766 59454 78818
rect 60386 78766 60398 78818
rect 60450 78766 60462 78818
rect 64306 78766 64318 78818
rect 64370 78766 64382 78818
rect 69570 78766 69582 78818
rect 69634 78766 69646 78818
rect 82002 78766 82014 78818
rect 82066 78766 82078 78818
rect 53342 78754 53394 78766
rect 62302 78754 62354 78766
rect 68574 78754 68626 78766
rect 75966 78754 76018 78766
rect 83022 78754 83074 78766
rect 83806 78818 83858 78830
rect 86718 78818 86770 78830
rect 93214 78818 93266 78830
rect 85698 78766 85710 78818
rect 85762 78766 85774 78818
rect 86146 78766 86158 78818
rect 86210 78766 86222 78818
rect 87490 78766 87502 78818
rect 87554 78766 87566 78818
rect 88386 78766 88398 78818
rect 88450 78766 88462 78818
rect 91634 78766 91646 78818
rect 91698 78766 91710 78818
rect 94882 78766 94894 78818
rect 94946 78766 94958 78818
rect 83806 78754 83858 78766
rect 86718 78754 86770 78766
rect 93214 78754 93266 78766
rect 49310 78706 49362 78718
rect 49310 78642 49362 78654
rect 50654 78706 50706 78718
rect 50654 78642 50706 78654
rect 50766 78706 50818 78718
rect 50766 78642 50818 78654
rect 51662 78706 51714 78718
rect 51662 78642 51714 78654
rect 53566 78706 53618 78718
rect 53566 78642 53618 78654
rect 53678 78706 53730 78718
rect 53678 78642 53730 78654
rect 58830 78706 58882 78718
rect 67790 78706 67842 78718
rect 65090 78654 65102 78706
rect 65154 78654 65166 78706
rect 58830 78642 58882 78654
rect 67790 78642 67842 78654
rect 67902 78706 67954 78718
rect 67902 78642 67954 78654
rect 75182 78706 75234 78718
rect 75182 78642 75234 78654
rect 75518 78706 75570 78718
rect 75518 78642 75570 78654
rect 76302 78706 76354 78718
rect 76302 78642 76354 78654
rect 83358 78706 83410 78718
rect 83358 78642 83410 78654
rect 84030 78706 84082 78718
rect 84030 78642 84082 78654
rect 84142 78706 84194 78718
rect 84142 78642 84194 78654
rect 91870 78706 91922 78718
rect 91870 78642 91922 78654
rect 49758 78594 49810 78606
rect 49758 78530 49810 78542
rect 50206 78594 50258 78606
rect 50206 78530 50258 78542
rect 50990 78594 51042 78606
rect 50990 78530 51042 78542
rect 51326 78594 51378 78606
rect 51326 78530 51378 78542
rect 51550 78594 51602 78606
rect 51550 78530 51602 78542
rect 52334 78594 52386 78606
rect 52334 78530 52386 78542
rect 54238 78594 54290 78606
rect 61294 78594 61346 78606
rect 58370 78542 58382 78594
rect 58434 78542 58446 78594
rect 54238 78530 54290 78542
rect 61294 78530 61346 78542
rect 61742 78594 61794 78606
rect 61742 78530 61794 78542
rect 62638 78594 62690 78606
rect 62638 78530 62690 78542
rect 68126 78594 68178 78606
rect 68126 78530 68178 78542
rect 76190 78594 76242 78606
rect 76190 78530 76242 78542
rect 83246 78594 83298 78606
rect 89518 78594 89570 78606
rect 86258 78542 86270 78594
rect 86322 78542 86334 78594
rect 83246 78530 83298 78542
rect 89518 78530 89570 78542
rect 93550 78594 93602 78606
rect 93550 78530 93602 78542
rect 1344 78426 98560 78460
rect 1344 78374 19838 78426
rect 19890 78374 19942 78426
rect 19994 78374 20046 78426
rect 20098 78374 50558 78426
rect 50610 78374 50662 78426
rect 50714 78374 50766 78426
rect 50818 78374 81278 78426
rect 81330 78374 81382 78426
rect 81434 78374 81486 78426
rect 81538 78374 98560 78426
rect 1344 78340 98560 78374
rect 48862 78258 48914 78270
rect 48862 78194 48914 78206
rect 49982 78258 50034 78270
rect 49982 78194 50034 78206
rect 50766 78258 50818 78270
rect 50766 78194 50818 78206
rect 53678 78258 53730 78270
rect 53678 78194 53730 78206
rect 54126 78258 54178 78270
rect 54126 78194 54178 78206
rect 63422 78258 63474 78270
rect 63422 78194 63474 78206
rect 65326 78258 65378 78270
rect 65326 78194 65378 78206
rect 66334 78258 66386 78270
rect 69806 78258 69858 78270
rect 67666 78206 67678 78258
rect 67730 78206 67742 78258
rect 66334 78194 66386 78206
rect 69806 78194 69858 78206
rect 70030 78258 70082 78270
rect 70030 78194 70082 78206
rect 70590 78258 70642 78270
rect 70590 78194 70642 78206
rect 96350 78258 96402 78270
rect 96350 78194 96402 78206
rect 48302 78146 48354 78158
rect 48302 78082 48354 78094
rect 49646 78146 49698 78158
rect 49646 78082 49698 78094
rect 49758 78146 49810 78158
rect 49758 78082 49810 78094
rect 50430 78146 50482 78158
rect 50430 78082 50482 78094
rect 50542 78146 50594 78158
rect 50542 78082 50594 78094
rect 51326 78146 51378 78158
rect 51326 78082 51378 78094
rect 52110 78146 52162 78158
rect 52110 78082 52162 78094
rect 54910 78146 54962 78158
rect 54910 78082 54962 78094
rect 56590 78146 56642 78158
rect 56590 78082 56642 78094
rect 58046 78146 58098 78158
rect 58046 78082 58098 78094
rect 59278 78146 59330 78158
rect 65550 78146 65602 78158
rect 60274 78094 60286 78146
rect 60338 78094 60350 78146
rect 59278 78082 59330 78094
rect 65550 78082 65602 78094
rect 69022 78146 69074 78158
rect 69022 78082 69074 78094
rect 69358 78146 69410 78158
rect 69358 78082 69410 78094
rect 70142 78146 70194 78158
rect 70142 78082 70194 78094
rect 77310 78146 77362 78158
rect 89406 78146 89458 78158
rect 78306 78094 78318 78146
rect 78370 78094 78382 78146
rect 77310 78082 77362 78094
rect 89406 78082 89458 78094
rect 89518 78146 89570 78158
rect 93538 78094 93550 78146
rect 93602 78094 93614 78146
rect 95442 78094 95454 78146
rect 95506 78094 95518 78146
rect 89518 78082 89570 78094
rect 51214 78034 51266 78046
rect 51214 77970 51266 77982
rect 51550 78034 51602 78046
rect 51550 77970 51602 77982
rect 51886 78034 51938 78046
rect 51886 77970 51938 77982
rect 52222 78034 52274 78046
rect 52222 77970 52274 77982
rect 52670 78034 52722 78046
rect 52670 77970 52722 77982
rect 55022 78034 55074 78046
rect 55022 77970 55074 77982
rect 56366 78034 56418 78046
rect 56366 77970 56418 77982
rect 56702 78034 56754 78046
rect 56702 77970 56754 77982
rect 57822 78034 57874 78046
rect 57822 77970 57874 77982
rect 58158 78034 58210 78046
rect 60958 78034 61010 78046
rect 65662 78034 65714 78046
rect 59714 77982 59726 78034
rect 59778 77982 59790 78034
rect 60050 77982 60062 78034
rect 60114 77982 60126 78034
rect 61506 77982 61518 78034
rect 61570 77982 61582 78034
rect 62290 77982 62302 78034
rect 62354 77982 62366 78034
rect 58158 77970 58210 77982
rect 60958 77970 61010 77982
rect 65662 77970 65714 77982
rect 66110 78034 66162 78046
rect 66110 77970 66162 77982
rect 66446 78034 66498 78046
rect 66446 77970 66498 77982
rect 66894 78034 66946 78046
rect 66894 77970 66946 77982
rect 68014 78034 68066 78046
rect 68014 77970 68066 77982
rect 68462 78034 68514 78046
rect 68462 77970 68514 77982
rect 71598 78034 71650 78046
rect 78766 78034 78818 78046
rect 89182 78034 89234 78046
rect 72034 77982 72046 78034
rect 72098 77982 72110 78034
rect 73938 77982 73950 78034
rect 74002 77982 74014 78034
rect 77746 77982 77758 78034
rect 77810 77982 77822 78034
rect 78082 77982 78094 78034
rect 78146 77982 78158 78034
rect 79314 77982 79326 78034
rect 79378 77982 79390 78034
rect 80322 77982 80334 78034
rect 80386 77982 80398 78034
rect 81442 77982 81454 78034
rect 81506 77982 81518 78034
rect 87602 77982 87614 78034
rect 87666 77982 87678 78034
rect 88386 77982 88398 78034
rect 88450 77982 88462 78034
rect 94322 77982 94334 78034
rect 94386 77982 94398 78034
rect 95218 77982 95230 78034
rect 95282 77982 95294 78034
rect 71598 77970 71650 77982
rect 78766 77970 78818 77982
rect 89182 77970 89234 77982
rect 53118 77922 53170 77934
rect 53118 77858 53170 77870
rect 57374 77922 57426 77934
rect 57374 77858 57426 77870
rect 58606 77922 58658 77934
rect 58606 77858 58658 77870
rect 62974 77922 63026 77934
rect 62974 77858 63026 77870
rect 71038 77922 71090 77934
rect 71038 77858 71090 77870
rect 73278 77922 73330 77934
rect 84702 77922 84754 77934
rect 74610 77870 74622 77922
rect 74674 77870 74686 77922
rect 76738 77870 76750 77922
rect 76802 77870 76814 77922
rect 82114 77870 82126 77922
rect 82178 77870 82190 77922
rect 84242 77870 84254 77922
rect 84306 77870 84318 77922
rect 85474 77870 85486 77922
rect 85538 77870 85550 77922
rect 91410 77870 91422 77922
rect 91474 77870 91486 77922
rect 73278 77858 73330 77870
rect 84702 77858 84754 77870
rect 54910 77810 54962 77822
rect 54910 77746 54962 77758
rect 96014 77810 96066 77822
rect 96014 77746 96066 77758
rect 1344 77642 98560 77676
rect 1344 77590 4478 77642
rect 4530 77590 4582 77642
rect 4634 77590 4686 77642
rect 4738 77590 35198 77642
rect 35250 77590 35302 77642
rect 35354 77590 35406 77642
rect 35458 77590 65918 77642
rect 65970 77590 66022 77642
rect 66074 77590 66126 77642
rect 66178 77590 96638 77642
rect 96690 77590 96742 77642
rect 96794 77590 96846 77642
rect 96898 77590 98560 77642
rect 1344 77556 98560 77590
rect 72830 77474 72882 77486
rect 57474 77422 57486 77474
rect 57538 77471 57550 77474
rect 58258 77471 58270 77474
rect 57538 77425 58270 77471
rect 57538 77422 57550 77425
rect 58258 77422 58270 77425
rect 58322 77422 58334 77474
rect 94322 77422 94334 77474
rect 94386 77471 94398 77474
rect 94882 77471 94894 77474
rect 94386 77425 94894 77471
rect 94386 77422 94398 77425
rect 94882 77422 94894 77425
rect 94946 77422 94958 77474
rect 72830 77410 72882 77422
rect 69246 77362 69298 77374
rect 52658 77310 52670 77362
rect 52722 77310 52734 77362
rect 55122 77310 55134 77362
rect 55186 77310 55198 77362
rect 57250 77310 57262 77362
rect 57314 77310 57326 77362
rect 69246 77298 69298 77310
rect 79886 77362 79938 77374
rect 79886 77298 79938 77310
rect 82238 77362 82290 77374
rect 88734 77362 88786 77374
rect 85250 77310 85262 77362
rect 85314 77310 85326 77362
rect 82238 77298 82290 77310
rect 88734 77298 88786 77310
rect 94670 77362 94722 77374
rect 94670 77298 94722 77310
rect 57710 77250 57762 77262
rect 49858 77198 49870 77250
rect 49922 77198 49934 77250
rect 54338 77198 54350 77250
rect 54402 77198 54414 77250
rect 57710 77186 57762 77198
rect 62078 77250 62130 77262
rect 70814 77250 70866 77262
rect 67890 77198 67902 77250
rect 67954 77198 67966 77250
rect 62078 77186 62130 77198
rect 70814 77186 70866 77198
rect 71822 77250 71874 77262
rect 71822 77186 71874 77198
rect 76526 77250 76578 77262
rect 76526 77186 76578 77198
rect 78878 77250 78930 77262
rect 78878 77186 78930 77198
rect 80446 77250 80498 77262
rect 80446 77186 80498 77198
rect 80782 77250 80834 77262
rect 80782 77186 80834 77198
rect 84366 77250 84418 77262
rect 88162 77198 88174 77250
rect 88226 77198 88238 77250
rect 93314 77198 93326 77250
rect 93378 77198 93390 77250
rect 84366 77186 84418 77198
rect 72158 77138 72210 77150
rect 50530 77086 50542 77138
rect 50594 77086 50606 77138
rect 64306 77086 64318 77138
rect 64370 77086 64382 77138
rect 72158 77074 72210 77086
rect 72718 77138 72770 77150
rect 72718 77074 72770 77086
rect 72830 77138 72882 77150
rect 72830 77074 72882 77086
rect 74958 77138 75010 77150
rect 74958 77074 75010 77086
rect 75518 77138 75570 77150
rect 75518 77074 75570 77086
rect 77198 77138 77250 77150
rect 77198 77074 77250 77086
rect 77534 77138 77586 77150
rect 77534 77074 77586 77086
rect 77982 77138 78034 77150
rect 77982 77074 78034 77086
rect 78206 77138 78258 77150
rect 78206 77074 78258 77086
rect 78318 77138 78370 77150
rect 81454 77138 81506 77150
rect 79202 77086 79214 77138
rect 79266 77086 79278 77138
rect 78318 77074 78370 77086
rect 81454 77074 81506 77086
rect 81790 77138 81842 77150
rect 81790 77074 81842 77086
rect 83022 77138 83074 77150
rect 83022 77074 83074 77086
rect 83134 77138 83186 77150
rect 87378 77086 87390 77138
rect 87442 77086 87454 77138
rect 83134 77074 83186 77086
rect 53342 77026 53394 77038
rect 53342 76962 53394 76974
rect 53790 77026 53842 77038
rect 53790 76962 53842 76974
rect 58158 77026 58210 77038
rect 58158 76962 58210 76974
rect 58606 77026 58658 77038
rect 58606 76962 58658 76974
rect 68350 77026 68402 77038
rect 68350 76962 68402 76974
rect 69694 77026 69746 77038
rect 69694 76962 69746 76974
rect 71262 77026 71314 77038
rect 71262 76962 71314 76974
rect 71934 77026 71986 77038
rect 71934 76962 71986 76974
rect 74286 77026 74338 77038
rect 74286 76962 74338 76974
rect 74622 77026 74674 77038
rect 74622 76962 74674 76974
rect 74846 77026 74898 77038
rect 74846 76962 74898 76974
rect 75854 77026 75906 77038
rect 75854 76962 75906 76974
rect 77422 77026 77474 77038
rect 77422 76962 77474 76974
rect 81678 77026 81730 77038
rect 81678 76962 81730 76974
rect 83358 77026 83410 77038
rect 83358 76962 83410 76974
rect 84030 77026 84082 77038
rect 84030 76962 84082 76974
rect 84254 77026 84306 77038
rect 84254 76962 84306 76974
rect 90862 77026 90914 77038
rect 90862 76962 90914 76974
rect 92542 77026 92594 77038
rect 92542 76962 92594 76974
rect 93550 77026 93602 77038
rect 93550 76962 93602 76974
rect 95006 77026 95058 77038
rect 95006 76962 95058 76974
rect 1344 76858 98560 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 81278 76858
rect 81330 76806 81382 76858
rect 81434 76806 81486 76858
rect 81538 76806 98560 76858
rect 1344 76772 98560 76806
rect 58382 76690 58434 76702
rect 58382 76626 58434 76638
rect 58942 76690 58994 76702
rect 58942 76626 58994 76638
rect 63534 76690 63586 76702
rect 63534 76626 63586 76638
rect 64542 76690 64594 76702
rect 64542 76626 64594 76638
rect 65438 76690 65490 76702
rect 65438 76626 65490 76638
rect 67006 76690 67058 76702
rect 67006 76626 67058 76638
rect 76974 76690 77026 76702
rect 76974 76626 77026 76638
rect 77758 76690 77810 76702
rect 77758 76626 77810 76638
rect 78542 76690 78594 76702
rect 78542 76626 78594 76638
rect 80222 76690 80274 76702
rect 80222 76626 80274 76638
rect 87278 76690 87330 76702
rect 87278 76626 87330 76638
rect 87614 76690 87666 76702
rect 87614 76626 87666 76638
rect 57598 76578 57650 76590
rect 57598 76514 57650 76526
rect 57710 76578 57762 76590
rect 57710 76514 57762 76526
rect 64766 76578 64818 76590
rect 64766 76514 64818 76526
rect 66446 76578 66498 76590
rect 66446 76514 66498 76526
rect 66558 76578 66610 76590
rect 66558 76514 66610 76526
rect 67230 76578 67282 76590
rect 81454 76578 81506 76590
rect 74386 76526 74398 76578
rect 74450 76526 74462 76578
rect 67230 76514 67282 76526
rect 81454 76514 81506 76526
rect 82238 76578 82290 76590
rect 82238 76514 82290 76526
rect 82798 76578 82850 76590
rect 87054 76578 87106 76590
rect 84242 76526 84254 76578
rect 84306 76526 84318 76578
rect 82798 76514 82850 76526
rect 87054 76514 87106 76526
rect 90302 76578 90354 76590
rect 90302 76514 90354 76526
rect 58494 76466 58546 76478
rect 52882 76414 52894 76466
rect 52946 76414 52958 76466
rect 58494 76402 58546 76414
rect 64430 76466 64482 76478
rect 64430 76402 64482 76414
rect 65774 76466 65826 76478
rect 65774 76402 65826 76414
rect 67342 76466 67394 76478
rect 71598 76466 71650 76478
rect 81230 76466 81282 76478
rect 68114 76414 68126 76466
rect 68178 76414 68190 76466
rect 73714 76414 73726 76466
rect 73778 76414 73790 76466
rect 67342 76402 67394 76414
rect 71598 76402 71650 76414
rect 81230 76402 81282 76414
rect 81566 76466 81618 76478
rect 81566 76402 81618 76414
rect 82350 76466 82402 76478
rect 86942 76466 86994 76478
rect 83570 76414 83582 76466
rect 83634 76414 83646 76466
rect 82350 76402 82402 76414
rect 86942 76402 86994 76414
rect 90638 76466 90690 76478
rect 91858 76414 91870 76466
rect 91922 76414 91934 76466
rect 90638 76402 90690 76414
rect 50878 76354 50930 76366
rect 63870 76354 63922 76366
rect 72158 76354 72210 76366
rect 56466 76302 56478 76354
rect 56530 76302 56542 76354
rect 68898 76302 68910 76354
rect 68962 76302 68974 76354
rect 71026 76302 71038 76354
rect 71090 76302 71102 76354
rect 50878 76290 50930 76302
rect 63870 76290 63922 76302
rect 72158 76290 72210 76302
rect 72606 76354 72658 76366
rect 80558 76354 80610 76366
rect 97134 76354 97186 76366
rect 76514 76302 76526 76354
rect 76578 76302 76590 76354
rect 86370 76302 86382 76354
rect 86434 76302 86446 76354
rect 94882 76302 94894 76354
rect 94946 76302 94958 76354
rect 72606 76290 72658 76302
rect 80558 76290 80610 76302
rect 97134 76290 97186 76302
rect 57598 76242 57650 76254
rect 57598 76178 57650 76190
rect 58382 76242 58434 76254
rect 58382 76178 58434 76190
rect 66446 76242 66498 76254
rect 66446 76178 66498 76190
rect 82238 76242 82290 76254
rect 82238 76178 82290 76190
rect 1344 76074 98560 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 96638 76074
rect 96690 76022 96742 76074
rect 96794 76022 96846 76074
rect 96898 76022 98560 76074
rect 1344 75988 98560 76022
rect 97134 75906 97186 75918
rect 67554 75854 67566 75906
rect 67618 75903 67630 75906
rect 68114 75903 68126 75906
rect 67618 75857 68126 75903
rect 67618 75854 67630 75857
rect 68114 75854 68126 75857
rect 68178 75854 68190 75906
rect 97134 75842 97186 75854
rect 62974 75794 63026 75806
rect 67566 75794 67618 75806
rect 50530 75742 50542 75794
rect 50594 75742 50606 75794
rect 52658 75742 52670 75794
rect 52722 75742 52734 75794
rect 56690 75742 56702 75794
rect 56754 75742 56766 75794
rect 58034 75742 58046 75794
rect 58098 75742 58110 75794
rect 60162 75742 60174 75794
rect 60226 75742 60238 75794
rect 64530 75742 64542 75794
rect 64594 75742 64606 75794
rect 66658 75742 66670 75794
rect 66722 75742 66734 75794
rect 62974 75730 63026 75742
rect 67566 75730 67618 75742
rect 70142 75794 70194 75806
rect 70142 75730 70194 75742
rect 70590 75794 70642 75806
rect 70590 75730 70642 75742
rect 71262 75794 71314 75806
rect 71262 75730 71314 75742
rect 73390 75794 73442 75806
rect 73390 75730 73442 75742
rect 73726 75794 73778 75806
rect 86718 75794 86770 75806
rect 79762 75742 79774 75794
rect 79826 75742 79838 75794
rect 81890 75742 81902 75794
rect 81954 75742 81966 75794
rect 90290 75742 90302 75794
rect 90354 75742 90366 75794
rect 92418 75742 92430 75794
rect 92482 75742 92494 75794
rect 93202 75742 93214 75794
rect 93266 75742 93278 75794
rect 95330 75742 95342 75794
rect 95394 75742 95406 75794
rect 73726 75730 73778 75742
rect 86718 75730 86770 75742
rect 67118 75682 67170 75694
rect 49858 75630 49870 75682
rect 49922 75630 49934 75682
rect 53778 75630 53790 75682
rect 53842 75630 53854 75682
rect 57362 75630 57374 75682
rect 57426 75630 57438 75682
rect 63746 75630 63758 75682
rect 63810 75630 63822 75682
rect 67118 75618 67170 75630
rect 68014 75682 68066 75694
rect 68014 75618 68066 75630
rect 74622 75682 74674 75694
rect 74622 75618 74674 75630
rect 76302 75682 76354 75694
rect 82350 75682 82402 75694
rect 79090 75630 79102 75682
rect 79154 75630 79166 75682
rect 76302 75618 76354 75630
rect 82350 75618 82402 75630
rect 82686 75682 82738 75694
rect 82686 75618 82738 75630
rect 83470 75682 83522 75694
rect 83470 75618 83522 75630
rect 84590 75682 84642 75694
rect 84590 75618 84642 75630
rect 85598 75682 85650 75694
rect 85598 75618 85650 75630
rect 86046 75682 86098 75694
rect 86046 75618 86098 75630
rect 86382 75682 86434 75694
rect 89506 75630 89518 75682
rect 89570 75630 89582 75682
rect 96002 75630 96014 75682
rect 96066 75630 96078 75682
rect 86382 75618 86434 75630
rect 62526 75570 62578 75582
rect 54562 75518 54574 75570
rect 54626 75518 54638 75570
rect 62526 75506 62578 75518
rect 69358 75570 69410 75582
rect 69358 75506 69410 75518
rect 69694 75570 69746 75582
rect 69694 75506 69746 75518
rect 74286 75570 74338 75582
rect 74286 75506 74338 75518
rect 75070 75570 75122 75582
rect 75070 75506 75122 75518
rect 75406 75570 75458 75582
rect 75406 75506 75458 75518
rect 75966 75570 76018 75582
rect 75966 75506 76018 75518
rect 76078 75570 76130 75582
rect 76078 75506 76130 75518
rect 84254 75570 84306 75582
rect 84254 75506 84306 75518
rect 85262 75570 85314 75582
rect 85262 75506 85314 75518
rect 85374 75570 85426 75582
rect 85374 75506 85426 75518
rect 86158 75570 86210 75582
rect 97346 75518 97358 75570
rect 97410 75518 97422 75570
rect 97794 75518 97806 75570
rect 97858 75518 97870 75570
rect 86158 75506 86210 75518
rect 62190 75458 62242 75470
rect 62190 75394 62242 75406
rect 74398 75458 74450 75470
rect 74398 75394 74450 75406
rect 82574 75458 82626 75470
rect 82574 75394 82626 75406
rect 83134 75458 83186 75470
rect 83134 75394 83186 75406
rect 83358 75458 83410 75470
rect 83358 75394 83410 75406
rect 84366 75458 84418 75470
rect 84366 75394 84418 75406
rect 89070 75458 89122 75470
rect 89070 75394 89122 75406
rect 96798 75458 96850 75470
rect 96798 75394 96850 75406
rect 1344 75290 98560 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 81278 75290
rect 81330 75238 81382 75290
rect 81434 75238 81486 75290
rect 81538 75238 98560 75290
rect 1344 75204 98560 75238
rect 53342 75122 53394 75134
rect 53342 75058 53394 75070
rect 53566 75122 53618 75134
rect 53566 75058 53618 75070
rect 54126 75122 54178 75134
rect 54126 75058 54178 75070
rect 54910 75122 54962 75134
rect 54910 75058 54962 75070
rect 55134 75122 55186 75134
rect 55134 75058 55186 75070
rect 55694 75122 55746 75134
rect 55694 75058 55746 75070
rect 57374 75122 57426 75134
rect 57374 75058 57426 75070
rect 57822 75122 57874 75134
rect 57822 75058 57874 75070
rect 65438 75122 65490 75134
rect 65438 75058 65490 75070
rect 66222 75122 66274 75134
rect 66222 75058 66274 75070
rect 70590 75122 70642 75134
rect 70590 75058 70642 75070
rect 74622 75122 74674 75134
rect 74622 75058 74674 75070
rect 76078 75122 76130 75134
rect 76078 75058 76130 75070
rect 85150 75122 85202 75134
rect 85150 75058 85202 75070
rect 91422 75122 91474 75134
rect 91422 75058 91474 75070
rect 93438 75122 93490 75134
rect 93438 75058 93490 75070
rect 54350 75010 54402 75022
rect 50754 74958 50766 75010
rect 50818 74958 50830 75010
rect 54350 74946 54402 74958
rect 55918 75010 55970 75022
rect 55918 74946 55970 74958
rect 56030 75010 56082 75022
rect 56030 74946 56082 74958
rect 65774 75010 65826 75022
rect 75070 75010 75122 75022
rect 71474 74958 71486 75010
rect 71538 74958 71550 75010
rect 65774 74946 65826 74958
rect 75070 74946 75122 74958
rect 88510 75010 88562 75022
rect 95566 75010 95618 75022
rect 89954 74958 89966 75010
rect 90018 74958 90030 75010
rect 90514 74958 90526 75010
rect 90578 74958 90590 75010
rect 91970 74958 91982 75010
rect 92034 74958 92046 75010
rect 92306 74958 92318 75010
rect 92370 74958 92382 75010
rect 93986 74958 93998 75010
rect 94050 74958 94062 75010
rect 94322 74958 94334 75010
rect 94386 74958 94398 75010
rect 88510 74946 88562 74958
rect 95566 74946 95618 74958
rect 95902 75010 95954 75022
rect 95902 74946 95954 74958
rect 53678 74898 53730 74910
rect 49970 74846 49982 74898
rect 50034 74846 50046 74898
rect 53678 74834 53730 74846
rect 54462 74898 54514 74910
rect 54462 74834 54514 74846
rect 55246 74898 55298 74910
rect 64318 74898 64370 74910
rect 70926 74898 70978 74910
rect 74286 74898 74338 74910
rect 89406 74898 89458 74910
rect 60610 74846 60622 74898
rect 60674 74846 60686 74898
rect 66994 74846 67006 74898
rect 67058 74846 67070 74898
rect 71698 74846 71710 74898
rect 71762 74846 71774 74898
rect 81778 74846 81790 74898
rect 81842 74846 81854 74898
rect 88274 74846 88286 74898
rect 88338 74846 88350 74898
rect 55246 74834 55298 74846
rect 64318 74834 64370 74846
rect 70926 74834 70978 74846
rect 74286 74834 74338 74846
rect 89406 74834 89458 74846
rect 56478 74786 56530 74798
rect 63982 74786 64034 74798
rect 72270 74786 72322 74798
rect 52882 74734 52894 74786
rect 52946 74734 52958 74786
rect 61282 74734 61294 74786
rect 61346 74734 61358 74786
rect 63410 74734 63422 74786
rect 63474 74734 63486 74786
rect 67778 74734 67790 74786
rect 67842 74734 67854 74786
rect 69906 74734 69918 74786
rect 69970 74734 69982 74786
rect 56478 74722 56530 74734
rect 63982 74722 64034 74734
rect 72270 74722 72322 74734
rect 73726 74786 73778 74798
rect 73726 74722 73778 74734
rect 75742 74786 75794 74798
rect 75742 74722 75794 74734
rect 81342 74786 81394 74798
rect 89742 74786 89794 74798
rect 82562 74734 82574 74786
rect 82626 74734 82638 74786
rect 84690 74734 84702 74786
rect 84754 74734 84766 74786
rect 81342 74722 81394 74734
rect 89742 74722 89794 74734
rect 96350 74786 96402 74798
rect 96350 74722 96402 74734
rect 97134 74786 97186 74798
rect 97134 74722 97186 74734
rect 91758 74674 91810 74686
rect 91758 74610 91810 74622
rect 93774 74674 93826 74686
rect 93774 74610 93826 74622
rect 1344 74506 98560 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 96638 74506
rect 96690 74454 96742 74506
rect 96794 74454 96846 74506
rect 96898 74454 98560 74506
rect 1344 74420 98560 74454
rect 82562 74286 82574 74338
rect 82626 74335 82638 74338
rect 82898 74335 82910 74338
rect 82626 74289 82910 74335
rect 82626 74286 82638 74289
rect 82898 74286 82910 74289
rect 82962 74286 82974 74338
rect 50206 74226 50258 74238
rect 50206 74162 50258 74174
rect 53342 74226 53394 74238
rect 53342 74162 53394 74174
rect 53902 74226 53954 74238
rect 53902 74162 53954 74174
rect 54350 74226 54402 74238
rect 54350 74162 54402 74174
rect 54798 74226 54850 74238
rect 82238 74226 82290 74238
rect 67554 74174 67566 74226
rect 67618 74174 67630 74226
rect 54798 74162 54850 74174
rect 82238 74162 82290 74174
rect 82686 74226 82738 74238
rect 82686 74162 82738 74174
rect 84366 74226 84418 74238
rect 91646 74226 91698 74238
rect 88610 74174 88622 74226
rect 88674 74174 88686 74226
rect 90738 74174 90750 74226
rect 90802 74174 90814 74226
rect 84366 74162 84418 74174
rect 91646 74162 91698 74174
rect 92094 74226 92146 74238
rect 92094 74162 92146 74174
rect 93102 74226 93154 74238
rect 93102 74162 93154 74174
rect 93550 74226 93602 74238
rect 95666 74174 95678 74226
rect 95730 74174 95742 74226
rect 97794 74174 97806 74226
rect 97858 74174 97870 74226
rect 93550 74162 93602 74174
rect 50654 74114 50706 74126
rect 50654 74050 50706 74062
rect 51326 74114 51378 74126
rect 51326 74050 51378 74062
rect 51662 74114 51714 74126
rect 51662 74050 51714 74062
rect 52110 74114 52162 74126
rect 52110 74050 52162 74062
rect 52446 74114 52498 74126
rect 61518 74114 61570 74126
rect 60386 74062 60398 74114
rect 60450 74062 60462 74114
rect 52446 74050 52498 74062
rect 61518 74050 61570 74062
rect 61854 74114 61906 74126
rect 69806 74114 69858 74126
rect 76526 74114 76578 74126
rect 62402 74062 62414 74114
rect 62466 74062 62478 74114
rect 63858 74062 63870 74114
rect 63922 74062 63934 74114
rect 74834 74062 74846 74114
rect 74898 74062 74910 74114
rect 76066 74062 76078 74114
rect 76130 74062 76142 74114
rect 61854 74050 61906 74062
rect 69806 74050 69858 74062
rect 76526 74050 76578 74062
rect 83022 74114 83074 74126
rect 83022 74050 83074 74062
rect 83358 74114 83410 74126
rect 87826 74062 87838 74114
rect 87890 74062 87902 74114
rect 94882 74062 94894 74114
rect 94946 74062 94958 74114
rect 83358 74050 83410 74062
rect 50990 74002 51042 74014
rect 50990 73938 51042 73950
rect 59726 74002 59778 74014
rect 59726 73938 59778 73950
rect 60622 74002 60674 74014
rect 69470 74002 69522 74014
rect 71934 74002 71986 74014
rect 62626 73950 62638 74002
rect 62690 73950 62702 74002
rect 70018 73950 70030 74002
rect 70082 73950 70094 74002
rect 70578 73950 70590 74002
rect 70642 73950 70654 74002
rect 60622 73938 60674 73950
rect 69470 73938 69522 73950
rect 71934 73938 71986 73950
rect 72270 74002 72322 74014
rect 72270 73938 72322 73950
rect 72718 74002 72770 74014
rect 72718 73938 72770 73950
rect 77422 74002 77474 74014
rect 77422 73938 77474 73950
rect 78542 74002 78594 74014
rect 78542 73938 78594 73950
rect 83806 74002 83858 74014
rect 83806 73938 83858 73950
rect 91310 74002 91362 74014
rect 91310 73938 91362 73950
rect 50766 73890 50818 73902
rect 50766 73826 50818 73838
rect 51550 73890 51602 73902
rect 51550 73826 51602 73838
rect 52334 73890 52386 73902
rect 52334 73826 52386 73838
rect 71262 73890 71314 73902
rect 71262 73826 71314 73838
rect 75070 73890 75122 73902
rect 75070 73826 75122 73838
rect 78206 73890 78258 73902
rect 78206 73826 78258 73838
rect 83246 73890 83298 73902
rect 83246 73826 83298 73838
rect 93998 73890 94050 73902
rect 93998 73826 94050 73838
rect 1344 73722 98560 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 81278 73722
rect 81330 73670 81382 73722
rect 81434 73670 81486 73722
rect 81538 73670 98560 73722
rect 1344 73636 98560 73670
rect 58270 73554 58322 73566
rect 58270 73490 58322 73502
rect 59502 73554 59554 73566
rect 59502 73490 59554 73502
rect 65326 73554 65378 73566
rect 65326 73490 65378 73502
rect 68238 73554 68290 73566
rect 68238 73490 68290 73502
rect 79326 73554 79378 73566
rect 79326 73490 79378 73502
rect 91086 73554 91138 73566
rect 91086 73490 91138 73502
rect 56030 73442 56082 73454
rect 68574 73442 68626 73454
rect 81790 73442 81842 73454
rect 62178 73390 62190 73442
rect 62242 73390 62254 73442
rect 75058 73390 75070 73442
rect 75122 73390 75134 73442
rect 78306 73390 78318 73442
rect 78370 73390 78382 73442
rect 78754 73390 78766 73442
rect 78818 73390 78830 73442
rect 56030 73378 56082 73390
rect 68574 73378 68626 73390
rect 81790 73378 81842 73390
rect 83246 73442 83298 73454
rect 83246 73378 83298 73390
rect 88174 73442 88226 73454
rect 91982 73442 92034 73454
rect 89954 73390 89966 73442
rect 90018 73390 90030 73442
rect 90514 73390 90526 73442
rect 90578 73390 90590 73442
rect 88174 73378 88226 73390
rect 91982 73378 92034 73390
rect 93662 73442 93714 73454
rect 97246 73442 97298 73454
rect 95778 73390 95790 73442
rect 95842 73390 95854 73442
rect 96338 73390 96350 73442
rect 96402 73390 96414 73442
rect 93662 73378 93714 73390
rect 97246 73378 97298 73390
rect 56366 73330 56418 73342
rect 73726 73330 73778 73342
rect 88510 73330 88562 73342
rect 61506 73278 61518 73330
rect 61570 73278 61582 73330
rect 74386 73278 74398 73330
rect 74450 73278 74462 73330
rect 81554 73278 81566 73330
rect 81618 73278 81630 73330
rect 83010 73278 83022 73330
rect 83074 73278 83086 73330
rect 56366 73266 56418 73278
rect 73726 73266 73778 73278
rect 88510 73266 88562 73278
rect 89406 73330 89458 73342
rect 95230 73330 95282 73342
rect 91746 73278 91758 73330
rect 91810 73278 91822 73330
rect 89406 73266 89458 73278
rect 95230 73266 95282 73278
rect 97582 73330 97634 73342
rect 97582 73266 97634 73278
rect 51326 73218 51378 73230
rect 51326 73154 51378 73166
rect 51886 73218 51938 73230
rect 51886 73154 51938 73166
rect 57486 73218 57538 73230
rect 57486 73154 57538 73166
rect 57822 73218 57874 73230
rect 57822 73154 57874 73166
rect 60846 73218 60898 73230
rect 71150 73218 71202 73230
rect 64306 73166 64318 73218
rect 64370 73166 64382 73218
rect 60846 73154 60898 73166
rect 71150 73154 71202 73166
rect 72494 73218 72546 73230
rect 72494 73154 72546 73166
rect 73390 73218 73442 73230
rect 79998 73218 80050 73230
rect 77186 73166 77198 73218
rect 77250 73166 77262 73218
rect 73390 73154 73442 73166
rect 79998 73154 80050 73166
rect 94222 73218 94274 73230
rect 94222 73154 94274 73166
rect 94670 73218 94722 73230
rect 94670 73154 94722 73166
rect 78990 73106 79042 73118
rect 78990 73042 79042 73054
rect 89742 73106 89794 73118
rect 95566 73106 95618 73118
rect 94210 73054 94222 73106
rect 94274 73103 94286 73106
rect 94882 73103 94894 73106
rect 94274 73057 94894 73103
rect 94274 73054 94286 73057
rect 94882 73054 94894 73057
rect 94946 73054 94958 73106
rect 89742 73042 89794 73054
rect 95566 73042 95618 73054
rect 1344 72938 98560 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 96638 72938
rect 96690 72886 96742 72938
rect 96794 72886 96846 72938
rect 96898 72886 98560 72938
rect 1344 72852 98560 72886
rect 58046 72770 58098 72782
rect 58046 72706 58098 72718
rect 62078 72770 62130 72782
rect 62078 72706 62130 72718
rect 64766 72770 64818 72782
rect 64766 72706 64818 72718
rect 74846 72770 74898 72782
rect 74846 72706 74898 72718
rect 59726 72658 59778 72670
rect 59726 72594 59778 72606
rect 71710 72658 71762 72670
rect 77870 72658 77922 72670
rect 73490 72606 73502 72658
rect 73554 72606 73566 72658
rect 94882 72606 94894 72658
rect 94946 72606 94958 72658
rect 97010 72606 97022 72658
rect 97074 72606 97086 72658
rect 71710 72594 71762 72606
rect 77870 72594 77922 72606
rect 56478 72546 56530 72558
rect 58382 72546 58434 72558
rect 61742 72546 61794 72558
rect 64430 72546 64482 72558
rect 49746 72494 49758 72546
rect 49810 72494 49822 72546
rect 57138 72494 57150 72546
rect 57202 72494 57214 72546
rect 59154 72494 59166 72546
rect 59218 72494 59230 72546
rect 60386 72494 60398 72546
rect 60450 72494 60462 72546
rect 62738 72494 62750 72546
rect 62802 72494 62814 72546
rect 56478 72482 56530 72494
rect 58382 72482 58434 72494
rect 61742 72482 61794 72494
rect 64430 72482 64482 72494
rect 72270 72546 72322 72558
rect 72270 72482 72322 72494
rect 73950 72546 74002 72558
rect 73950 72482 74002 72494
rect 75182 72546 75234 72558
rect 75618 72494 75630 72546
rect 75682 72494 75694 72546
rect 83906 72494 83918 72546
rect 83970 72494 83982 72546
rect 87154 72494 87166 72546
rect 87218 72494 87230 72546
rect 97682 72494 97694 72546
rect 97746 72494 97758 72546
rect 75182 72482 75234 72494
rect 55470 72434 55522 72446
rect 55470 72370 55522 72382
rect 56142 72434 56194 72446
rect 70814 72434 70866 72446
rect 57250 72382 57262 72434
rect 57314 72382 57326 72434
rect 59042 72382 59054 72434
rect 59106 72382 59118 72434
rect 62850 72382 62862 72434
rect 62914 72382 62926 72434
rect 63634 72382 63646 72434
rect 63698 72382 63710 72434
rect 64194 72382 64206 72434
rect 64258 72382 64270 72434
rect 75954 72382 75966 72434
rect 76018 72382 76030 72434
rect 78978 72382 78990 72434
rect 79042 72382 79054 72434
rect 89170 72382 89182 72434
rect 89234 72382 89246 72434
rect 56142 72370 56194 72382
rect 70814 72370 70866 72382
rect 49982 72322 50034 72334
rect 49982 72258 50034 72270
rect 54686 72322 54738 72334
rect 54686 72258 54738 72270
rect 55134 72322 55186 72334
rect 55134 72258 55186 72270
rect 60622 72322 60674 72334
rect 60622 72258 60674 72270
rect 65326 72322 65378 72334
rect 65326 72258 65378 72270
rect 65774 72322 65826 72334
rect 65774 72258 65826 72270
rect 69246 72322 69298 72334
rect 69246 72258 69298 72270
rect 70478 72322 70530 72334
rect 70478 72258 70530 72270
rect 72830 72322 72882 72334
rect 72830 72258 72882 72270
rect 76526 72322 76578 72334
rect 76526 72258 76578 72270
rect 77198 72322 77250 72334
rect 77198 72258 77250 72270
rect 84478 72322 84530 72334
rect 84478 72258 84530 72270
rect 86606 72322 86658 72334
rect 86606 72258 86658 72270
rect 94110 72322 94162 72334
rect 94110 72258 94162 72270
rect 1344 72154 98560 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 81278 72154
rect 81330 72102 81382 72154
rect 81434 72102 81486 72154
rect 81538 72102 98560 72154
rect 1344 72068 98560 72102
rect 50430 71986 50482 71998
rect 50430 71922 50482 71934
rect 63646 71986 63698 71998
rect 63646 71922 63698 71934
rect 73838 71986 73890 71998
rect 73838 71922 73890 71934
rect 68910 71874 68962 71886
rect 51538 71822 51550 71874
rect 51602 71822 51614 71874
rect 54562 71822 54574 71874
rect 54626 71822 54638 71874
rect 70242 71822 70254 71874
rect 70306 71822 70318 71874
rect 78418 71822 78430 71874
rect 78482 71822 78494 71874
rect 82114 71822 82126 71874
rect 82178 71822 82190 71874
rect 92530 71822 92542 71874
rect 92594 71822 92606 71874
rect 68910 71810 68962 71822
rect 51426 71710 51438 71762
rect 51490 71710 51502 71762
rect 53778 71710 53790 71762
rect 53842 71710 53854 71762
rect 62738 71710 62750 71762
rect 62802 71710 62814 71762
rect 68674 71710 68686 71762
rect 68738 71710 68750 71762
rect 69570 71710 69582 71762
rect 69634 71710 69646 71762
rect 77634 71710 77646 71762
rect 77698 71710 77710 71762
rect 81330 71710 81342 71762
rect 81394 71710 81406 71762
rect 89842 71710 89854 71762
rect 89906 71710 89918 71762
rect 52110 71650 52162 71662
rect 52110 71586 52162 71598
rect 52670 71650 52722 71662
rect 52670 71586 52722 71598
rect 53342 71650 53394 71662
rect 63198 71650 63250 71662
rect 56690 71598 56702 71650
rect 56754 71598 56766 71650
rect 58818 71598 58830 71650
rect 58882 71598 58894 71650
rect 53342 71586 53394 71598
rect 63198 71586 63250 71598
rect 66110 71650 66162 71662
rect 66110 71586 66162 71598
rect 68014 71650 68066 71662
rect 73278 71650 73330 71662
rect 74846 71650 74898 71662
rect 72370 71598 72382 71650
rect 72434 71598 72446 71650
rect 74274 71598 74286 71650
rect 74338 71598 74350 71650
rect 68014 71586 68066 71598
rect 73278 71586 73330 71598
rect 74846 71586 74898 71598
rect 75294 71650 75346 71662
rect 75294 71586 75346 71598
rect 75742 71650 75794 71662
rect 75742 71586 75794 71598
rect 76302 71650 76354 71662
rect 76302 71586 76354 71598
rect 76638 71650 76690 71662
rect 95566 71650 95618 71662
rect 80546 71598 80558 71650
rect 80610 71598 80622 71650
rect 84242 71598 84254 71650
rect 84306 71598 84318 71650
rect 76638 71586 76690 71598
rect 95566 71586 95618 71598
rect 50766 71538 50818 71550
rect 74834 71486 74846 71538
rect 74898 71535 74910 71538
rect 75282 71535 75294 71538
rect 74898 71489 75294 71535
rect 74898 71486 74910 71489
rect 75282 71486 75294 71489
rect 75346 71535 75358 71538
rect 76738 71535 76750 71538
rect 75346 71489 76750 71535
rect 75346 71486 75358 71489
rect 76738 71486 76750 71489
rect 76802 71486 76814 71538
rect 50766 71474 50818 71486
rect 1344 71370 98560 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 96638 71370
rect 96690 71318 96742 71370
rect 96794 71318 96846 71370
rect 96898 71318 98560 71370
rect 1344 71284 98560 71318
rect 82014 71202 82066 71214
rect 82014 71138 82066 71150
rect 82350 71202 82402 71214
rect 82350 71138 82402 71150
rect 85374 71202 85426 71214
rect 85374 71138 85426 71150
rect 85710 71202 85762 71214
rect 85710 71138 85762 71150
rect 92318 71202 92370 71214
rect 92318 71138 92370 71150
rect 67230 71090 67282 71102
rect 77198 71090 77250 71102
rect 51650 71038 51662 71090
rect 51714 71038 51726 71090
rect 55794 71038 55806 71090
rect 55858 71038 55870 71090
rect 57922 71038 57934 71090
rect 57986 71038 57998 71090
rect 62178 71038 62190 71090
rect 62242 71038 62254 71090
rect 64306 71038 64318 71090
rect 64370 71038 64382 71090
rect 71362 71038 71374 71090
rect 71426 71038 71438 71090
rect 67230 71026 67282 71038
rect 77198 71026 77250 71038
rect 80334 71090 80386 71102
rect 80334 71026 80386 71038
rect 80782 71090 80834 71102
rect 93662 71090 93714 71102
rect 88386 71038 88398 71090
rect 88450 71038 88462 71090
rect 90514 71038 90526 71090
rect 90578 71038 90590 71090
rect 80782 71026 80834 71038
rect 93662 71026 93714 71038
rect 93998 71090 94050 71102
rect 93998 71026 94050 71038
rect 96462 71090 96514 71102
rect 96462 71026 96514 71038
rect 58942 70978 58994 70990
rect 76078 70978 76130 70990
rect 91982 70978 92034 70990
rect 48850 70926 48862 70978
rect 48914 70926 48926 70978
rect 55122 70926 55134 70978
rect 55186 70926 55198 70978
rect 61506 70926 61518 70978
rect 61570 70926 61582 70978
rect 69346 70926 69358 70978
rect 69410 70926 69422 70978
rect 75282 70926 75294 70978
rect 75346 70926 75358 70978
rect 83010 70926 83022 70978
rect 83074 70926 83086 70978
rect 87714 70926 87726 70978
rect 87778 70926 87790 70978
rect 91298 70926 91310 70978
rect 91362 70926 91374 70978
rect 58942 70914 58994 70926
rect 76078 70914 76130 70926
rect 91982 70914 92034 70926
rect 93102 70978 93154 70990
rect 93102 70914 93154 70926
rect 47854 70866 47906 70878
rect 47854 70802 47906 70814
rect 48190 70866 48242 70878
rect 53566 70866 53618 70878
rect 49522 70814 49534 70866
rect 49586 70814 49598 70866
rect 48190 70802 48242 70814
rect 53566 70802 53618 70814
rect 53902 70866 53954 70878
rect 65662 70866 65714 70878
rect 59154 70814 59166 70866
rect 59218 70814 59230 70866
rect 59490 70814 59502 70866
rect 59554 70814 59566 70866
rect 53902 70802 53954 70814
rect 65662 70802 65714 70814
rect 66334 70866 66386 70878
rect 66334 70802 66386 70814
rect 66670 70866 66722 70878
rect 66670 70802 66722 70814
rect 68238 70866 68290 70878
rect 68238 70802 68290 70814
rect 68574 70866 68626 70878
rect 94782 70866 94834 70878
rect 82898 70814 82910 70866
rect 82962 70814 82974 70866
rect 85922 70814 85934 70866
rect 85986 70814 85998 70866
rect 86258 70814 86270 70866
rect 86322 70814 86334 70866
rect 91186 70814 91198 70866
rect 91250 70814 91262 70866
rect 68574 70802 68626 70814
rect 94782 70802 94834 70814
rect 95118 70866 95170 70878
rect 95118 70802 95170 70814
rect 95678 70866 95730 70878
rect 95678 70802 95730 70814
rect 52110 70754 52162 70766
rect 52110 70690 52162 70702
rect 52670 70754 52722 70766
rect 52670 70690 52722 70702
rect 58606 70754 58658 70766
rect 58606 70690 58658 70702
rect 60286 70754 60338 70766
rect 60286 70690 60338 70702
rect 64766 70754 64818 70766
rect 64766 70690 64818 70702
rect 65326 70754 65378 70766
rect 65326 70690 65378 70702
rect 67790 70754 67842 70766
rect 67790 70690 67842 70702
rect 75518 70754 75570 70766
rect 75518 70690 75570 70702
rect 76414 70754 76466 70766
rect 76414 70690 76466 70702
rect 77758 70754 77810 70766
rect 77758 70690 77810 70702
rect 81454 70754 81506 70766
rect 81454 70690 81506 70702
rect 83694 70754 83746 70766
rect 83694 70690 83746 70702
rect 84590 70754 84642 70766
rect 84590 70690 84642 70702
rect 87054 70754 87106 70766
rect 87054 70690 87106 70702
rect 96014 70754 96066 70766
rect 96014 70690 96066 70702
rect 1344 70586 98560 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 81278 70586
rect 81330 70534 81382 70586
rect 81434 70534 81486 70586
rect 81538 70534 98560 70586
rect 1344 70500 98560 70534
rect 63870 70418 63922 70430
rect 63870 70354 63922 70366
rect 66222 70418 66274 70430
rect 66222 70354 66274 70366
rect 71486 70418 71538 70430
rect 71486 70354 71538 70366
rect 72606 70418 72658 70430
rect 72606 70354 72658 70366
rect 81230 70418 81282 70430
rect 81230 70354 81282 70366
rect 88062 70418 88114 70430
rect 88062 70354 88114 70366
rect 89294 70418 89346 70430
rect 89294 70354 89346 70366
rect 94782 70418 94834 70430
rect 94782 70354 94834 70366
rect 90302 70306 90354 70318
rect 56466 70254 56478 70306
rect 56530 70254 56542 70306
rect 58482 70254 58494 70306
rect 58546 70254 58558 70306
rect 66770 70254 66782 70306
rect 66834 70254 66846 70306
rect 67330 70254 67342 70306
rect 67394 70254 67406 70306
rect 68898 70254 68910 70306
rect 68962 70254 68974 70306
rect 76178 70254 76190 70306
rect 76242 70254 76254 70306
rect 83234 70254 83246 70306
rect 83298 70254 83310 70306
rect 93090 70254 93102 70306
rect 93154 70254 93166 70306
rect 95330 70254 95342 70306
rect 95394 70254 95406 70306
rect 95666 70254 95678 70306
rect 95730 70254 95742 70306
rect 90302 70242 90354 70254
rect 59278 70194 59330 70206
rect 72046 70194 72098 70206
rect 87166 70194 87218 70206
rect 52882 70142 52894 70194
rect 52946 70142 52958 70194
rect 58706 70142 58718 70194
rect 58770 70142 58782 70194
rect 60610 70142 60622 70194
rect 60674 70142 60686 70194
rect 68114 70142 68126 70194
rect 68178 70142 68190 70194
rect 76962 70142 76974 70194
rect 77026 70142 77038 70194
rect 77634 70142 77646 70194
rect 77698 70142 77710 70194
rect 82562 70142 82574 70194
rect 82626 70142 82638 70194
rect 59278 70130 59330 70142
rect 72046 70130 72098 70142
rect 87166 70130 87218 70142
rect 89630 70194 89682 70206
rect 89630 70130 89682 70142
rect 90190 70194 90242 70206
rect 90190 70130 90242 70142
rect 90526 70194 90578 70206
rect 96462 70194 96514 70206
rect 93874 70142 93886 70194
rect 93938 70142 93950 70194
rect 90526 70130 90578 70142
rect 96462 70130 96514 70142
rect 59726 70082 59778 70094
rect 73390 70082 73442 70094
rect 87726 70082 87778 70094
rect 61282 70030 61294 70082
rect 61346 70030 61358 70082
rect 63410 70030 63422 70082
rect 63474 70030 63486 70082
rect 71026 70030 71038 70082
rect 71090 70030 71102 70082
rect 74050 70030 74062 70082
rect 74114 70030 74126 70082
rect 78306 70030 78318 70082
rect 78370 70030 78382 70082
rect 80434 70030 80446 70082
rect 80498 70030 80510 70082
rect 85362 70030 85374 70082
rect 85426 70030 85438 70082
rect 59726 70018 59778 70030
rect 73390 70018 73442 70030
rect 87726 70018 87778 70030
rect 88510 70082 88562 70094
rect 95118 70082 95170 70094
rect 90962 70030 90974 70082
rect 91026 70030 91038 70082
rect 88510 70018 88562 70030
rect 95118 70018 95170 70030
rect 97134 70082 97186 70094
rect 97134 70018 97186 70030
rect 57598 69970 57650 69982
rect 57598 69906 57650 69918
rect 57934 69970 57986 69982
rect 66558 69970 66610 69982
rect 59042 69918 59054 69970
rect 59106 69967 59118 69970
rect 59826 69967 59838 69970
rect 59106 69921 59838 69967
rect 59106 69918 59118 69921
rect 59826 69918 59838 69921
rect 59890 69918 59902 69970
rect 57934 69906 57986 69918
rect 66558 69906 66610 69918
rect 1344 69802 98560 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 96638 69802
rect 96690 69750 96742 69802
rect 96794 69750 96846 69802
rect 96898 69750 98560 69802
rect 1344 69716 98560 69750
rect 70254 69634 70306 69646
rect 70254 69570 70306 69582
rect 72158 69634 72210 69646
rect 72158 69570 72210 69582
rect 72494 69634 72546 69646
rect 72494 69570 72546 69582
rect 75742 69634 75794 69646
rect 75742 69570 75794 69582
rect 84366 69634 84418 69646
rect 84366 69570 84418 69582
rect 60398 69522 60450 69534
rect 69246 69522 69298 69534
rect 52434 69470 52446 69522
rect 52498 69470 52510 69522
rect 56466 69470 56478 69522
rect 56530 69470 56542 69522
rect 59938 69470 59950 69522
rect 60002 69470 60014 69522
rect 63858 69470 63870 69522
rect 63922 69470 63934 69522
rect 60398 69458 60450 69470
rect 69246 69458 69298 69470
rect 81230 69522 81282 69534
rect 81230 69458 81282 69470
rect 82686 69522 82738 69534
rect 94110 69522 94162 69534
rect 86034 69470 86046 69522
rect 86098 69470 86110 69522
rect 88162 69470 88174 69522
rect 88226 69470 88238 69522
rect 89506 69470 89518 69522
rect 89570 69470 89582 69522
rect 94882 69470 94894 69522
rect 94946 69470 94958 69522
rect 97010 69470 97022 69522
rect 97074 69470 97086 69522
rect 82686 69458 82738 69470
rect 94110 69458 94162 69470
rect 70590 69410 70642 69422
rect 75406 69410 75458 69422
rect 49522 69358 49534 69410
rect 49586 69358 49598 69410
rect 53666 69358 53678 69410
rect 53730 69358 53742 69410
rect 57138 69358 57150 69410
rect 57202 69358 57214 69410
rect 65426 69358 65438 69410
rect 65490 69358 65502 69410
rect 71250 69358 71262 69410
rect 71314 69358 71326 69410
rect 73266 69358 73278 69410
rect 73330 69358 73342 69410
rect 70590 69346 70642 69358
rect 75406 69346 75458 69358
rect 78206 69410 78258 69422
rect 78206 69346 78258 69358
rect 79102 69410 79154 69422
rect 84478 69410 84530 69422
rect 89070 69410 89122 69422
rect 81890 69358 81902 69410
rect 81954 69358 81966 69410
rect 85250 69358 85262 69410
rect 85314 69358 85326 69410
rect 92418 69358 92430 69410
rect 92482 69358 92494 69410
rect 93426 69358 93438 69410
rect 93490 69358 93502 69410
rect 97682 69358 97694 69410
rect 97746 69358 97758 69410
rect 79102 69346 79154 69358
rect 84478 69346 84530 69358
rect 89070 69346 89122 69358
rect 67566 69298 67618 69310
rect 50306 69246 50318 69298
rect 50370 69246 50382 69298
rect 54338 69246 54350 69298
rect 54402 69246 54414 69298
rect 57810 69246 57822 69298
rect 57874 69246 57886 69298
rect 67566 69234 67618 69246
rect 67678 69298 67730 69310
rect 67678 69234 67730 69246
rect 68574 69298 68626 69310
rect 82126 69298 82178 69310
rect 71362 69246 71374 69298
rect 71426 69246 71438 69298
rect 73042 69246 73054 69298
rect 73106 69246 73118 69298
rect 74834 69246 74846 69298
rect 74898 69246 74910 69298
rect 75170 69246 75182 69298
rect 75234 69246 75246 69298
rect 77410 69246 77422 69298
rect 77474 69246 77486 69298
rect 77970 69246 77982 69298
rect 78034 69246 78046 69298
rect 68574 69234 68626 69246
rect 82126 69234 82178 69246
rect 83246 69298 83298 69310
rect 83246 69234 83298 69246
rect 83358 69298 83410 69310
rect 83358 69234 83410 69246
rect 88734 69298 88786 69310
rect 88734 69234 88786 69246
rect 88846 69298 88898 69310
rect 93214 69298 93266 69310
rect 91634 69246 91646 69298
rect 91698 69246 91710 69298
rect 88846 69234 88898 69246
rect 93214 69234 93266 69246
rect 67902 69186 67954 69198
rect 67902 69122 67954 69134
rect 68238 69186 68290 69198
rect 68238 69122 68290 69134
rect 68462 69186 68514 69198
rect 68462 69122 68514 69134
rect 73950 69186 74002 69198
rect 73950 69122 74002 69134
rect 76302 69186 76354 69198
rect 76302 69122 76354 69134
rect 78542 69186 78594 69198
rect 78542 69122 78594 69134
rect 79550 69186 79602 69198
rect 79550 69122 79602 69134
rect 79998 69186 80050 69198
rect 79998 69122 80050 69134
rect 83582 69186 83634 69198
rect 83582 69122 83634 69134
rect 84366 69186 84418 69198
rect 84366 69122 84418 69134
rect 1344 69018 98560 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 81278 69018
rect 81330 68966 81382 69018
rect 81434 68966 81486 69018
rect 81538 68966 98560 69018
rect 1344 68932 98560 68966
rect 50206 68850 50258 68862
rect 50206 68786 50258 68798
rect 52670 68850 52722 68862
rect 52670 68786 52722 68798
rect 53678 68850 53730 68862
rect 53678 68786 53730 68798
rect 54238 68850 54290 68862
rect 54238 68786 54290 68798
rect 55134 68850 55186 68862
rect 55134 68786 55186 68798
rect 56478 68850 56530 68862
rect 56478 68786 56530 68798
rect 57374 68850 57426 68862
rect 57374 68786 57426 68798
rect 60622 68850 60674 68862
rect 60622 68786 60674 68798
rect 61182 68850 61234 68862
rect 61182 68786 61234 68798
rect 65550 68850 65602 68862
rect 65550 68786 65602 68798
rect 73726 68850 73778 68862
rect 73726 68786 73778 68798
rect 74846 68850 74898 68862
rect 74846 68786 74898 68798
rect 77198 68850 77250 68862
rect 77198 68786 77250 68798
rect 90526 68850 90578 68862
rect 90526 68786 90578 68798
rect 52110 68738 52162 68750
rect 51314 68686 51326 68738
rect 51378 68686 51390 68738
rect 52110 68674 52162 68686
rect 54574 68738 54626 68750
rect 75742 68738 75794 68750
rect 63298 68686 63310 68738
rect 63362 68686 63374 68738
rect 54574 68674 54626 68686
rect 75742 68674 75794 68686
rect 78094 68738 78146 68750
rect 78094 68674 78146 68686
rect 79214 68738 79266 68750
rect 79214 68674 79266 68686
rect 79998 68738 80050 68750
rect 89618 68686 89630 68738
rect 89682 68686 89694 68738
rect 96226 68686 96238 68738
rect 96290 68686 96302 68738
rect 79998 68674 80050 68686
rect 51886 68626 51938 68638
rect 51202 68574 51214 68626
rect 51266 68574 51278 68626
rect 51886 68562 51938 68574
rect 52222 68626 52274 68638
rect 61518 68626 61570 68638
rect 55346 68574 55358 68626
rect 55410 68574 55422 68626
rect 56242 68574 56254 68626
rect 56306 68574 56318 68626
rect 52222 68562 52274 68574
rect 61518 68562 61570 68574
rect 62190 68626 62242 68638
rect 63870 68626 63922 68638
rect 74286 68626 74338 68638
rect 63186 68574 63198 68626
rect 63250 68574 63262 68626
rect 66098 68574 66110 68626
rect 66162 68574 66174 68626
rect 62190 68562 62242 68574
rect 63870 68562 63922 68574
rect 74286 68562 74338 68574
rect 75182 68626 75234 68638
rect 75182 68562 75234 68574
rect 76302 68626 76354 68638
rect 77758 68626 77810 68638
rect 76962 68574 76974 68626
rect 77026 68574 77038 68626
rect 76302 68562 76354 68574
rect 77758 68562 77810 68574
rect 79102 68626 79154 68638
rect 79102 68562 79154 68574
rect 79438 68626 79490 68638
rect 79438 68562 79490 68574
rect 79886 68626 79938 68638
rect 90190 68626 90242 68638
rect 87378 68574 87390 68626
rect 87442 68574 87454 68626
rect 89394 68574 89406 68626
rect 89458 68574 89470 68626
rect 91186 68574 91198 68626
rect 91250 68574 91262 68626
rect 79886 68562 79938 68574
rect 90190 68562 90242 68574
rect 53118 68514 53170 68526
rect 53118 68450 53170 68462
rect 64318 68514 64370 68526
rect 69582 68514 69634 68526
rect 66882 68462 66894 68514
rect 66946 68462 66958 68514
rect 69010 68462 69022 68514
rect 69074 68462 69086 68514
rect 64318 68450 64370 68462
rect 69582 68450 69634 68462
rect 69918 68514 69970 68526
rect 69918 68450 69970 68462
rect 70590 68514 70642 68526
rect 70590 68450 70642 68462
rect 71038 68514 71090 68526
rect 71038 68450 71090 68462
rect 71374 68514 71426 68526
rect 71374 68450 71426 68462
rect 71934 68514 71986 68526
rect 71934 68450 71986 68462
rect 72494 68514 72546 68526
rect 72494 68450 72546 68462
rect 78654 68514 78706 68526
rect 83458 68462 83470 68514
rect 83522 68462 83534 68514
rect 78654 68450 78706 68462
rect 50542 68402 50594 68414
rect 62526 68402 62578 68414
rect 52434 68350 52446 68402
rect 52498 68399 52510 68402
rect 52994 68399 53006 68402
rect 52498 68353 53006 68399
rect 52498 68350 52510 68353
rect 52994 68350 53006 68353
rect 53058 68350 53070 68402
rect 50542 68338 50594 68350
rect 62526 68338 62578 68350
rect 79998 68402 80050 68414
rect 79998 68338 80050 68350
rect 1344 68234 98560 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 96638 68234
rect 96690 68182 96742 68234
rect 96794 68182 96846 68234
rect 96898 68182 98560 68234
rect 1344 68148 98560 68182
rect 61854 68066 61906 68078
rect 52098 68014 52110 68066
rect 52162 68063 52174 68066
rect 52546 68063 52558 68066
rect 52162 68017 52558 68063
rect 52162 68014 52174 68017
rect 52546 68014 52558 68017
rect 52610 68014 52622 68066
rect 61854 68002 61906 68014
rect 68462 68066 68514 68078
rect 68462 68002 68514 68014
rect 59390 67954 59442 67966
rect 49634 67902 49646 67954
rect 49698 67902 49710 67954
rect 51762 67902 51774 67954
rect 51826 67902 51838 67954
rect 59390 67890 59442 67902
rect 63198 67954 63250 67966
rect 69246 67954 69298 67966
rect 73390 67954 73442 67966
rect 64866 67902 64878 67954
rect 64930 67902 64942 67954
rect 66994 67902 67006 67954
rect 67058 67902 67070 67954
rect 72594 67902 72606 67954
rect 72658 67902 72670 67954
rect 63198 67890 63250 67902
rect 69246 67890 69298 67902
rect 73390 67890 73442 67902
rect 75742 67954 75794 67966
rect 75742 67890 75794 67902
rect 76190 67954 76242 67966
rect 92094 67954 92146 67966
rect 77522 67902 77534 67954
rect 77586 67902 77598 67954
rect 88162 67902 88174 67954
rect 88226 67902 88238 67954
rect 88722 67902 88734 67954
rect 88786 67902 88798 67954
rect 90850 67902 90862 67954
rect 90914 67902 90926 67954
rect 93538 67902 93550 67954
rect 93602 67902 93614 67954
rect 95666 67902 95678 67954
rect 95730 67902 95742 67954
rect 76190 67890 76242 67902
rect 92094 67890 92146 67902
rect 67454 67842 67506 67854
rect 48962 67790 48974 67842
rect 49026 67790 49038 67842
rect 62290 67790 62302 67842
rect 62354 67790 62366 67842
rect 64082 67790 64094 67842
rect 64146 67790 64158 67842
rect 67454 67778 67506 67790
rect 67790 67842 67842 67854
rect 83022 67842 83074 67854
rect 72482 67790 72494 67842
rect 72546 67790 72558 67842
rect 73826 67790 73838 67842
rect 73890 67790 73902 67842
rect 82562 67790 82574 67842
rect 82626 67790 82638 67842
rect 67790 67778 67842 67790
rect 83022 67778 83074 67790
rect 84254 67842 84306 67854
rect 97358 67842 97410 67854
rect 85250 67790 85262 67842
rect 85314 67790 85326 67842
rect 91522 67790 91534 67842
rect 91586 67790 91598 67842
rect 96338 67790 96350 67842
rect 96402 67790 96414 67842
rect 84254 67778 84306 67790
rect 97358 67778 97410 67790
rect 60622 67730 60674 67742
rect 60622 67666 60674 67678
rect 61518 67730 61570 67742
rect 67678 67730 67730 67742
rect 62626 67678 62638 67730
rect 62690 67678 62702 67730
rect 61518 67666 61570 67678
rect 67678 67666 67730 67678
rect 68462 67730 68514 67742
rect 68462 67666 68514 67678
rect 68574 67730 68626 67742
rect 68574 67666 68626 67678
rect 72830 67730 72882 67742
rect 72830 67666 72882 67678
rect 83582 67730 83634 67742
rect 83582 67666 83634 67678
rect 83694 67730 83746 67742
rect 86034 67678 86046 67730
rect 86098 67678 86110 67730
rect 83694 67666 83746 67678
rect 52222 67618 52274 67630
rect 52222 67554 52274 67566
rect 52670 67618 52722 67630
rect 52670 67554 52722 67566
rect 53342 67618 53394 67630
rect 53342 67554 53394 67566
rect 53790 67618 53842 67630
rect 53790 67554 53842 67566
rect 54798 67618 54850 67630
rect 54798 67554 54850 67566
rect 60286 67618 60338 67630
rect 60286 67554 60338 67566
rect 69918 67618 69970 67630
rect 69918 67554 69970 67566
rect 70590 67618 70642 67630
rect 70590 67554 70642 67566
rect 71150 67618 71202 67630
rect 71150 67554 71202 67566
rect 71598 67618 71650 67630
rect 71598 67554 71650 67566
rect 72046 67618 72098 67630
rect 72046 67554 72098 67566
rect 74510 67618 74562 67630
rect 74510 67554 74562 67566
rect 74958 67618 75010 67630
rect 74958 67554 75010 67566
rect 75406 67618 75458 67630
rect 75406 67554 75458 67566
rect 83918 67618 83970 67630
rect 83918 67554 83970 67566
rect 96910 67618 96962 67630
rect 96910 67554 96962 67566
rect 1344 67450 98560 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 81278 67450
rect 81330 67398 81382 67450
rect 81434 67398 81486 67450
rect 81538 67398 98560 67450
rect 1344 67364 98560 67398
rect 50318 67282 50370 67294
rect 50318 67218 50370 67230
rect 51998 67282 52050 67294
rect 51998 67218 52050 67230
rect 52558 67282 52610 67294
rect 52558 67218 52610 67230
rect 52782 67282 52834 67294
rect 52782 67218 52834 67230
rect 63534 67282 63586 67294
rect 63534 67218 63586 67230
rect 71822 67282 71874 67294
rect 74510 67282 74562 67294
rect 73378 67230 73390 67282
rect 73442 67230 73454 67282
rect 71822 67218 71874 67230
rect 74510 67218 74562 67230
rect 76078 67282 76130 67294
rect 76078 67218 76130 67230
rect 83806 67282 83858 67294
rect 83806 67218 83858 67230
rect 85374 67282 85426 67294
rect 85374 67218 85426 67230
rect 86494 67282 86546 67294
rect 86494 67218 86546 67230
rect 49758 67170 49810 67182
rect 49758 67106 49810 67118
rect 51102 67170 51154 67182
rect 51102 67106 51154 67118
rect 51214 67170 51266 67182
rect 51214 67106 51266 67118
rect 51886 67170 51938 67182
rect 51886 67106 51938 67118
rect 52894 67170 52946 67182
rect 52894 67106 52946 67118
rect 53790 67170 53842 67182
rect 53790 67106 53842 67118
rect 54238 67170 54290 67182
rect 63086 67170 63138 67182
rect 69918 67170 69970 67182
rect 60498 67118 60510 67170
rect 60562 67118 60574 67170
rect 67330 67118 67342 67170
rect 67394 67118 67406 67170
rect 54238 67106 54290 67118
rect 63086 67106 63138 67118
rect 69918 67106 69970 67118
rect 70142 67170 70194 67182
rect 70142 67106 70194 67118
rect 70254 67170 70306 67182
rect 70254 67106 70306 67118
rect 73950 67170 74002 67182
rect 73950 67106 74002 67118
rect 75966 67170 76018 67182
rect 75966 67106 76018 67118
rect 77086 67170 77138 67182
rect 77086 67106 77138 67118
rect 81230 67170 81282 67182
rect 81230 67106 81282 67118
rect 81454 67170 81506 67182
rect 81454 67106 81506 67118
rect 83246 67170 83298 67182
rect 83246 67106 83298 67118
rect 84254 67170 84306 67182
rect 84254 67106 84306 67118
rect 84702 67170 84754 67182
rect 84702 67106 84754 67118
rect 85150 67170 85202 67182
rect 85150 67106 85202 67118
rect 85486 67170 85538 67182
rect 85486 67106 85538 67118
rect 86718 67170 86770 67182
rect 86718 67106 86770 67118
rect 87726 67170 87778 67182
rect 96350 67170 96402 67182
rect 91522 67118 91534 67170
rect 91586 67118 91598 67170
rect 95330 67118 95342 67170
rect 95394 67118 95406 67170
rect 87726 67106 87778 67118
rect 96350 67106 96402 67118
rect 48862 67058 48914 67070
rect 48862 66994 48914 67006
rect 50094 67058 50146 67070
rect 50094 66994 50146 67006
rect 50430 67058 50482 67070
rect 50430 66994 50482 67006
rect 51438 67058 51490 67070
rect 51438 66994 51490 67006
rect 52222 67058 52274 67070
rect 72158 67058 72210 67070
rect 76750 67058 76802 67070
rect 81566 67058 81618 67070
rect 59826 67006 59838 67058
rect 59890 67006 59902 67058
rect 66546 67006 66558 67058
rect 66610 67006 66622 67058
rect 74722 67006 74734 67058
rect 74786 67006 74798 67058
rect 77634 67006 77646 67058
rect 77698 67006 77710 67058
rect 52222 66994 52274 67006
rect 72158 66994 72210 67006
rect 76750 66994 76802 67006
rect 81566 66994 81618 67006
rect 83134 67058 83186 67070
rect 83134 66994 83186 67006
rect 86382 67058 86434 67070
rect 86382 66994 86434 67006
rect 87838 67058 87890 67070
rect 93986 67006 93998 67058
rect 94050 67006 94062 67058
rect 95218 67006 95230 67058
rect 95282 67006 95294 67058
rect 87838 66994 87890 67006
rect 48302 66946 48354 66958
rect 48302 66882 48354 66894
rect 53454 66946 53506 66958
rect 53454 66882 53506 66894
rect 58718 66946 58770 66958
rect 58718 66882 58770 66894
rect 59054 66946 59106 66958
rect 70702 66946 70754 66958
rect 62626 66894 62638 66946
rect 62690 66894 62702 66946
rect 69458 66894 69470 66946
rect 69522 66894 69534 66946
rect 59054 66882 59106 66894
rect 70702 66882 70754 66894
rect 71150 66946 71202 66958
rect 71150 66882 71202 66894
rect 72718 66946 72770 66958
rect 72718 66882 72770 66894
rect 75406 66946 75458 66958
rect 82014 66946 82066 66958
rect 78418 66894 78430 66946
rect 78482 66894 78494 66946
rect 80546 66894 80558 66946
rect 80610 66894 80622 66946
rect 75406 66882 75458 66894
rect 82014 66882 82066 66894
rect 87054 66946 87106 66958
rect 87054 66882 87106 66894
rect 88286 66946 88338 66958
rect 88286 66882 88338 66894
rect 96014 66946 96066 66958
rect 96014 66882 96066 66894
rect 97134 66946 97186 66958
rect 97134 66882 97186 66894
rect 97582 66946 97634 66958
rect 97582 66882 97634 66894
rect 73726 66834 73778 66846
rect 73726 66770 73778 66782
rect 76078 66834 76130 66846
rect 76078 66770 76130 66782
rect 83246 66834 83298 66846
rect 83246 66770 83298 66782
rect 87726 66834 87778 66846
rect 87726 66770 87778 66782
rect 1344 66666 98560 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 96638 66666
rect 96690 66614 96742 66666
rect 96794 66614 96846 66666
rect 96898 66614 98560 66666
rect 1344 66580 98560 66614
rect 65998 66498 66050 66510
rect 65998 66434 66050 66446
rect 74062 66498 74114 66510
rect 74062 66434 74114 66446
rect 90862 66498 90914 66510
rect 90862 66434 90914 66446
rect 57038 66386 57090 66398
rect 56466 66334 56478 66386
rect 56530 66334 56542 66386
rect 57038 66322 57090 66334
rect 58270 66386 58322 66398
rect 58270 66322 58322 66334
rect 63310 66386 63362 66398
rect 63310 66322 63362 66334
rect 67790 66386 67842 66398
rect 81902 66386 81954 66398
rect 73042 66334 73054 66386
rect 73106 66334 73118 66386
rect 79314 66334 79326 66386
rect 79378 66334 79390 66386
rect 81442 66334 81454 66386
rect 81506 66334 81518 66386
rect 67790 66322 67842 66334
rect 81902 66322 81954 66334
rect 82350 66386 82402 66398
rect 82350 66322 82402 66334
rect 85150 66386 85202 66398
rect 91870 66386 91922 66398
rect 88050 66334 88062 66386
rect 88114 66334 88126 66386
rect 90178 66334 90190 66386
rect 90242 66334 90254 66386
rect 85150 66322 85202 66334
rect 91870 66322 91922 66334
rect 94110 66386 94162 66398
rect 98030 66386 98082 66398
rect 97570 66334 97582 66386
rect 97634 66334 97646 66386
rect 94110 66322 94162 66334
rect 98030 66322 98082 66334
rect 49534 66274 49586 66286
rect 49534 66210 49586 66222
rect 52558 66274 52610 66286
rect 58942 66274 58994 66286
rect 61630 66274 61682 66286
rect 53554 66222 53566 66274
rect 53618 66222 53630 66274
rect 60386 66222 60398 66274
rect 60450 66222 60462 66274
rect 52558 66210 52610 66222
rect 58942 66210 58994 66222
rect 61630 66210 61682 66222
rect 61966 66274 62018 66286
rect 67566 66274 67618 66286
rect 66546 66222 66558 66274
rect 66610 66222 66622 66274
rect 61966 66210 62018 66222
rect 67566 66210 67618 66222
rect 68574 66274 68626 66286
rect 68574 66210 68626 66222
rect 69358 66274 69410 66286
rect 75518 66274 75570 66286
rect 85822 66274 85874 66286
rect 74050 66222 74062 66274
rect 74114 66222 74126 66274
rect 77410 66222 77422 66274
rect 77474 66222 77486 66274
rect 78530 66222 78542 66274
rect 78594 66222 78606 66274
rect 87378 66222 87390 66274
rect 87442 66222 87454 66274
rect 94658 66222 94670 66274
rect 94722 66222 94734 66274
rect 69358 66210 69410 66222
rect 75518 66210 75570 66222
rect 85822 66210 85874 66222
rect 49198 66162 49250 66174
rect 49198 66098 49250 66110
rect 50094 66162 50146 66174
rect 50094 66098 50146 66110
rect 50206 66162 50258 66174
rect 50206 66098 50258 66110
rect 50990 66162 51042 66174
rect 50990 66098 51042 66110
rect 51662 66162 51714 66174
rect 51662 66098 51714 66110
rect 51774 66162 51826 66174
rect 58830 66162 58882 66174
rect 67902 66162 67954 66174
rect 54338 66110 54350 66162
rect 54402 66110 54414 66162
rect 62290 66110 62302 66162
rect 62354 66110 62366 66162
rect 62626 66110 62638 66162
rect 62690 66110 62702 66162
rect 66770 66110 66782 66162
rect 66834 66110 66846 66162
rect 51774 66098 51826 66110
rect 58830 66098 58882 66110
rect 67902 66098 67954 66110
rect 69694 66162 69746 66174
rect 69694 66098 69746 66110
rect 73726 66162 73778 66174
rect 73726 66098 73778 66110
rect 74622 66162 74674 66174
rect 74622 66098 74674 66110
rect 74958 66162 75010 66174
rect 74958 66098 75010 66110
rect 75854 66162 75906 66174
rect 75854 66098 75906 66110
rect 84254 66162 84306 66174
rect 84254 66098 84306 66110
rect 84366 66162 84418 66174
rect 84366 66098 84418 66110
rect 90974 66162 91026 66174
rect 90974 66098 91026 66110
rect 91422 66162 91474 66174
rect 91422 66098 91474 66110
rect 93214 66162 93266 66174
rect 93214 66098 93266 66110
rect 93550 66162 93602 66174
rect 95442 66110 95454 66162
rect 95506 66110 95518 66162
rect 93550 66098 93602 66110
rect 49310 66050 49362 66062
rect 49310 65986 49362 65998
rect 49870 66050 49922 66062
rect 49870 65986 49922 65998
rect 50654 66050 50706 66062
rect 50654 65986 50706 65998
rect 50878 66050 50930 66062
rect 50878 65986 50930 65998
rect 51438 66050 51490 66062
rect 51438 65986 51490 65998
rect 52222 66050 52274 66062
rect 52222 65986 52274 65998
rect 52446 66050 52498 66062
rect 52446 65986 52498 65998
rect 58606 66050 58658 66062
rect 58606 65986 58658 65998
rect 59502 66050 59554 66062
rect 59502 65986 59554 65998
rect 60622 66050 60674 66062
rect 60622 65986 60674 65998
rect 64990 66050 65042 66062
rect 64990 65986 65042 65998
rect 65662 66050 65714 66062
rect 65662 65986 65714 65998
rect 67678 66050 67730 66062
rect 67678 65986 67730 65998
rect 68014 66050 68066 66062
rect 68014 65986 68066 65998
rect 69470 66050 69522 66062
rect 69470 65986 69522 65998
rect 70478 66050 70530 66062
rect 70478 65986 70530 65998
rect 70926 66050 70978 66062
rect 70926 65986 70978 65998
rect 71262 66050 71314 66062
rect 71262 65986 71314 65998
rect 71710 66050 71762 66062
rect 71710 65986 71762 65998
rect 72606 66050 72658 66062
rect 72606 65986 72658 65998
rect 76302 66050 76354 66062
rect 76302 65986 76354 65998
rect 77646 66050 77698 66062
rect 77646 65986 77698 65998
rect 82798 66050 82850 66062
rect 82798 65986 82850 65998
rect 83582 66050 83634 66062
rect 83582 65986 83634 65998
rect 84030 66050 84082 66062
rect 84030 65986 84082 65998
rect 85934 66050 85986 66062
rect 85934 65986 85986 65998
rect 86158 66050 86210 66062
rect 86158 65986 86210 65998
rect 86494 66050 86546 66062
rect 86494 65986 86546 65998
rect 90862 66050 90914 66062
rect 90862 65986 90914 65998
rect 92542 66050 92594 66062
rect 92542 65986 92594 65998
rect 1344 65882 98560 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 81278 65882
rect 81330 65830 81382 65882
rect 81434 65830 81486 65882
rect 81538 65830 98560 65882
rect 1344 65796 98560 65830
rect 53790 65714 53842 65726
rect 53790 65650 53842 65662
rect 54014 65714 54066 65726
rect 54014 65650 54066 65662
rect 55246 65714 55298 65726
rect 55246 65650 55298 65662
rect 63310 65714 63362 65726
rect 79102 65714 79154 65726
rect 73490 65662 73502 65714
rect 73554 65662 73566 65714
rect 63310 65650 63362 65662
rect 79102 65650 79154 65662
rect 79774 65714 79826 65726
rect 79774 65650 79826 65662
rect 88062 65714 88114 65726
rect 88062 65650 88114 65662
rect 90190 65714 90242 65726
rect 90190 65650 90242 65662
rect 90862 65714 90914 65726
rect 90862 65650 90914 65662
rect 91310 65714 91362 65726
rect 91310 65650 91362 65662
rect 94558 65714 94610 65726
rect 94558 65650 94610 65662
rect 53118 65602 53170 65614
rect 50306 65550 50318 65602
rect 50370 65550 50382 65602
rect 53118 65538 53170 65550
rect 53230 65602 53282 65614
rect 53230 65538 53282 65550
rect 54126 65602 54178 65614
rect 54126 65538 54178 65550
rect 55022 65602 55074 65614
rect 55022 65538 55074 65550
rect 58606 65602 58658 65614
rect 58606 65538 58658 65550
rect 58718 65602 58770 65614
rect 64318 65602 64370 65614
rect 60722 65550 60734 65602
rect 60786 65550 60798 65602
rect 58718 65538 58770 65550
rect 64318 65538 64370 65550
rect 64654 65602 64706 65614
rect 73950 65602 74002 65614
rect 66322 65550 66334 65602
rect 66386 65550 66398 65602
rect 64654 65538 64706 65550
rect 73950 65538 74002 65550
rect 75966 65602 76018 65614
rect 75966 65538 76018 65550
rect 77758 65602 77810 65614
rect 77758 65538 77810 65550
rect 79662 65602 79714 65614
rect 79662 65538 79714 65550
rect 86718 65602 86770 65614
rect 86718 65538 86770 65550
rect 86830 65602 86882 65614
rect 86830 65538 86882 65550
rect 89406 65602 89458 65614
rect 89406 65538 89458 65550
rect 89518 65602 89570 65614
rect 89518 65538 89570 65550
rect 90302 65602 90354 65614
rect 96338 65550 96350 65602
rect 96402 65550 96414 65602
rect 90302 65538 90354 65550
rect 54574 65490 54626 65502
rect 49634 65438 49646 65490
rect 49698 65438 49710 65490
rect 54574 65426 54626 65438
rect 55358 65490 55410 65502
rect 55358 65426 55410 65438
rect 55806 65490 55858 65502
rect 55806 65426 55858 65438
rect 57598 65490 57650 65502
rect 57598 65426 57650 65438
rect 57822 65490 57874 65502
rect 57822 65426 57874 65438
rect 58158 65490 58210 65502
rect 58158 65426 58210 65438
rect 58942 65490 58994 65502
rect 71150 65490 71202 65502
rect 59938 65438 59950 65490
rect 60002 65438 60014 65490
rect 69234 65438 69246 65490
rect 69298 65438 69310 65490
rect 58942 65426 58994 65438
rect 71150 65426 71202 65438
rect 71598 65490 71650 65502
rect 78094 65490 78146 65502
rect 79998 65490 80050 65502
rect 88174 65490 88226 65502
rect 74946 65438 74958 65490
rect 75010 65438 75022 65490
rect 77186 65438 77198 65490
rect 77250 65438 77262 65490
rect 78866 65438 78878 65490
rect 78930 65438 78942 65490
rect 83234 65438 83246 65490
rect 83298 65438 83310 65490
rect 83906 65438 83918 65490
rect 83970 65438 83982 65490
rect 71598 65426 71650 65438
rect 78094 65426 78146 65438
rect 79998 65426 80050 65438
rect 88174 65426 88226 65438
rect 89182 65490 89234 65502
rect 89182 65426 89234 65438
rect 89966 65490 90018 65502
rect 94322 65438 94334 65490
rect 94386 65438 94398 65490
rect 96114 65438 96126 65490
rect 96178 65438 96190 65490
rect 89966 65426 90018 65438
rect 56702 65378 56754 65390
rect 52434 65326 52446 65378
rect 52498 65326 52510 65378
rect 56702 65314 56754 65326
rect 57934 65378 57986 65390
rect 57934 65314 57986 65326
rect 59278 65378 59330 65390
rect 72046 65378 72098 65390
rect 62850 65326 62862 65378
rect 62914 65326 62926 65378
rect 59278 65314 59330 65326
rect 72046 65314 72098 65326
rect 72718 65378 72770 65390
rect 72718 65314 72770 65326
rect 80334 65378 80386 65390
rect 80334 65314 80386 65326
rect 81230 65378 81282 65390
rect 81230 65314 81282 65326
rect 81790 65378 81842 65390
rect 81790 65314 81842 65326
rect 82238 65378 82290 65390
rect 82238 65314 82290 65326
rect 82686 65378 82738 65390
rect 87390 65378 87442 65390
rect 86034 65326 86046 65378
rect 86098 65326 86110 65378
rect 82686 65314 82738 65326
rect 87390 65314 87442 65326
rect 93774 65378 93826 65390
rect 93774 65314 93826 65326
rect 53118 65266 53170 65278
rect 86718 65266 86770 65278
rect 70914 65214 70926 65266
rect 70978 65263 70990 65266
rect 71474 65263 71486 65266
rect 70978 65217 71486 65263
rect 70978 65214 70990 65217
rect 71474 65214 71486 65217
rect 71538 65214 71550 65266
rect 71698 65214 71710 65266
rect 71762 65263 71774 65266
rect 71922 65263 71934 65266
rect 71762 65217 71934 65263
rect 71762 65214 71774 65217
rect 71922 65214 71934 65217
rect 71986 65214 71998 65266
rect 53118 65202 53170 65214
rect 86718 65202 86770 65214
rect 88062 65266 88114 65278
rect 88062 65202 88114 65214
rect 95230 65266 95282 65278
rect 95230 65202 95282 65214
rect 95566 65266 95618 65278
rect 95566 65202 95618 65214
rect 1344 65098 98560 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 96638 65098
rect 96690 65046 96742 65098
rect 96794 65046 96846 65098
rect 96898 65046 98560 65098
rect 1344 65012 98560 65046
rect 81554 64878 81566 64930
rect 81618 64927 81630 64930
rect 82226 64927 82238 64930
rect 81618 64881 82238 64927
rect 81618 64878 81630 64881
rect 82226 64878 82238 64881
rect 82290 64878 82302 64930
rect 54126 64818 54178 64830
rect 49522 64766 49534 64818
rect 49586 64766 49598 64818
rect 51650 64766 51662 64818
rect 51714 64766 51726 64818
rect 54126 64754 54178 64766
rect 54574 64818 54626 64830
rect 54574 64754 54626 64766
rect 55470 64818 55522 64830
rect 61294 64818 61346 64830
rect 56354 64766 56366 64818
rect 56418 64766 56430 64818
rect 55470 64754 55522 64766
rect 61294 64754 61346 64766
rect 61742 64818 61794 64830
rect 67790 64818 67842 64830
rect 64754 64766 64766 64818
rect 64818 64766 64830 64818
rect 66882 64766 66894 64818
rect 66946 64766 66958 64818
rect 61742 64754 61794 64766
rect 67790 64754 67842 64766
rect 68126 64818 68178 64830
rect 68126 64754 68178 64766
rect 72046 64818 72098 64830
rect 72046 64754 72098 64766
rect 81566 64818 81618 64830
rect 81566 64754 81618 64766
rect 81902 64818 81954 64830
rect 81902 64754 81954 64766
rect 87054 64818 87106 64830
rect 97694 64818 97746 64830
rect 88610 64766 88622 64818
rect 88674 64766 88686 64818
rect 90738 64766 90750 64818
rect 90802 64766 90814 64818
rect 94210 64766 94222 64818
rect 94274 64766 94286 64818
rect 87054 64754 87106 64766
rect 97694 64754 97746 64766
rect 52110 64706 52162 64718
rect 48850 64654 48862 64706
rect 48914 64654 48926 64706
rect 52110 64642 52162 64654
rect 53342 64706 53394 64718
rect 53342 64642 53394 64654
rect 53678 64706 53730 64718
rect 53678 64642 53730 64654
rect 58046 64706 58098 64718
rect 58046 64642 58098 64654
rect 59838 64706 59890 64718
rect 59838 64642 59890 64654
rect 60622 64706 60674 64718
rect 69694 64706 69746 64718
rect 64082 64654 64094 64706
rect 64146 64654 64158 64706
rect 60622 64642 60674 64654
rect 69694 64642 69746 64654
rect 70814 64706 70866 64718
rect 70814 64642 70866 64654
rect 71262 64706 71314 64718
rect 71262 64642 71314 64654
rect 71598 64706 71650 64718
rect 71598 64642 71650 64654
rect 74398 64706 74450 64718
rect 74398 64642 74450 64654
rect 76414 64706 76466 64718
rect 80782 64706 80834 64718
rect 79986 64654 79998 64706
rect 80050 64654 80062 64706
rect 76414 64642 76466 64654
rect 80782 64642 80834 64654
rect 83246 64706 83298 64718
rect 83246 64642 83298 64654
rect 84254 64706 84306 64718
rect 84254 64642 84306 64654
rect 85486 64706 85538 64718
rect 87938 64654 87950 64706
rect 88002 64654 88014 64706
rect 97122 64654 97134 64706
rect 97186 64654 97198 64706
rect 85486 64642 85538 64654
rect 52446 64594 52498 64606
rect 52446 64530 52498 64542
rect 56926 64594 56978 64606
rect 56926 64530 56978 64542
rect 57486 64594 57538 64606
rect 57486 64530 57538 64542
rect 57822 64594 57874 64606
rect 57822 64530 57874 64542
rect 59390 64594 59442 64606
rect 59390 64530 59442 64542
rect 60510 64594 60562 64606
rect 60510 64530 60562 64542
rect 68574 64594 68626 64606
rect 68574 64530 68626 64542
rect 69358 64594 69410 64606
rect 69358 64530 69410 64542
rect 70478 64594 70530 64606
rect 70478 64530 70530 64542
rect 71486 64594 71538 64606
rect 71486 64530 71538 64542
rect 73278 64594 73330 64606
rect 73278 64530 73330 64542
rect 75854 64594 75906 64606
rect 75854 64530 75906 64542
rect 78206 64594 78258 64606
rect 78206 64530 78258 64542
rect 78990 64594 79042 64606
rect 78990 64530 79042 64542
rect 80894 64594 80946 64606
rect 80894 64530 80946 64542
rect 84142 64594 84194 64606
rect 84142 64530 84194 64542
rect 85374 64594 85426 64606
rect 85374 64530 85426 64542
rect 86046 64594 86098 64606
rect 86046 64530 86098 64542
rect 86270 64594 86322 64606
rect 86270 64530 86322 64542
rect 86606 64594 86658 64606
rect 96338 64542 96350 64594
rect 96402 64542 96414 64594
rect 86606 64530 86658 64542
rect 52334 64482 52386 64494
rect 52334 64418 52386 64430
rect 53566 64482 53618 64494
rect 53566 64418 53618 64430
rect 55022 64482 55074 64494
rect 55022 64418 55074 64430
rect 56366 64482 56418 64494
rect 56366 64418 56418 64430
rect 56478 64482 56530 64494
rect 56478 64418 56530 64430
rect 56702 64482 56754 64494
rect 56702 64418 56754 64430
rect 57710 64482 57762 64494
rect 57710 64418 57762 64430
rect 58494 64482 58546 64494
rect 58494 64418 58546 64430
rect 58942 64482 58994 64494
rect 58942 64418 58994 64430
rect 60286 64482 60338 64494
rect 77198 64482 77250 64494
rect 74162 64430 74174 64482
rect 74226 64430 74238 64482
rect 60286 64418 60338 64430
rect 77198 64418 77250 64430
rect 77870 64482 77922 64494
rect 77870 64418 77922 64430
rect 79326 64482 79378 64494
rect 79326 64418 79378 64430
rect 80222 64482 80274 64494
rect 80222 64418 80274 64430
rect 81118 64482 81170 64494
rect 81118 64418 81170 64430
rect 82350 64482 82402 64494
rect 82350 64418 82402 64430
rect 82910 64482 82962 64494
rect 82910 64418 82962 64430
rect 83918 64482 83970 64494
rect 83918 64418 83970 64430
rect 85150 64482 85202 64494
rect 85150 64418 85202 64430
rect 86382 64482 86434 64494
rect 86382 64418 86434 64430
rect 91198 64482 91250 64494
rect 91198 64418 91250 64430
rect 93662 64482 93714 64494
rect 93662 64418 93714 64430
rect 1344 64314 98560 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 81278 64314
rect 81330 64262 81382 64314
rect 81434 64262 81486 64314
rect 81538 64262 98560 64314
rect 1344 64228 98560 64262
rect 61630 64146 61682 64158
rect 58482 64094 58494 64146
rect 58546 64094 58558 64146
rect 61630 64082 61682 64094
rect 66222 64146 66274 64158
rect 66222 64082 66274 64094
rect 70926 64146 70978 64158
rect 70926 64082 70978 64094
rect 72158 64146 72210 64158
rect 72158 64082 72210 64094
rect 72718 64146 72770 64158
rect 77646 64146 77698 64158
rect 74386 64094 74398 64146
rect 74450 64094 74462 64146
rect 72718 64082 72770 64094
rect 77646 64082 77698 64094
rect 78206 64146 78258 64158
rect 79886 64146 79938 64158
rect 79314 64094 79326 64146
rect 79378 64094 79390 64146
rect 78206 64082 78258 64094
rect 79886 64082 79938 64094
rect 81902 64146 81954 64158
rect 81902 64082 81954 64094
rect 82014 64146 82066 64158
rect 82014 64082 82066 64094
rect 82910 64146 82962 64158
rect 82910 64082 82962 64094
rect 83022 64146 83074 64158
rect 83022 64082 83074 64094
rect 83134 64146 83186 64158
rect 83134 64082 83186 64094
rect 85038 64146 85090 64158
rect 85038 64082 85090 64094
rect 87054 64146 87106 64158
rect 87054 64082 87106 64094
rect 87502 64146 87554 64158
rect 87502 64082 87554 64094
rect 88398 64146 88450 64158
rect 93438 64146 93490 64158
rect 90290 64094 90302 64146
rect 90354 64094 90366 64146
rect 88398 64082 88450 64094
rect 93438 64082 93490 64094
rect 94558 64146 94610 64158
rect 94558 64082 94610 64094
rect 57486 64034 57538 64046
rect 50306 63982 50318 64034
rect 50370 63982 50382 64034
rect 54450 63982 54462 64034
rect 54514 63982 54526 64034
rect 57486 63970 57538 63982
rect 66670 64034 66722 64046
rect 70590 64034 70642 64046
rect 67666 63982 67678 64034
rect 67730 63982 67742 64034
rect 66670 63970 66722 63982
rect 70590 63970 70642 63982
rect 72382 64034 72434 64046
rect 72382 63970 72434 63982
rect 73950 64034 74002 64046
rect 73950 63970 74002 63982
rect 75966 64034 76018 64046
rect 75966 63970 76018 63982
rect 77758 64034 77810 64046
rect 77758 63970 77810 63982
rect 78430 64034 78482 64046
rect 78430 63970 78482 63982
rect 80222 64034 80274 64046
rect 80222 63970 80274 63982
rect 84814 64034 84866 64046
rect 96114 63982 96126 64034
rect 96178 63982 96190 64034
rect 84814 63970 84866 63982
rect 52894 63922 52946 63934
rect 55134 63922 55186 63934
rect 59166 63922 59218 63934
rect 61182 63922 61234 63934
rect 68350 63922 68402 63934
rect 71374 63922 71426 63934
rect 49522 63870 49534 63922
rect 49586 63870 49598 63922
rect 53890 63870 53902 63922
rect 53954 63870 53966 63922
rect 54226 63870 54238 63922
rect 54290 63870 54302 63922
rect 55682 63870 55694 63922
rect 55746 63870 55758 63922
rect 56578 63870 56590 63922
rect 56642 63870 56654 63922
rect 57922 63870 57934 63922
rect 57986 63870 57998 63922
rect 58258 63870 58270 63922
rect 58322 63870 58334 63922
rect 59714 63870 59726 63922
rect 59778 63870 59790 63922
rect 60498 63870 60510 63922
rect 60562 63870 60574 63922
rect 66994 63870 67006 63922
rect 67058 63870 67070 63922
rect 67442 63870 67454 63922
rect 67506 63870 67518 63922
rect 68786 63870 68798 63922
rect 68850 63870 68862 63922
rect 69682 63870 69694 63922
rect 69746 63870 69758 63922
rect 52894 63858 52946 63870
rect 55134 63858 55186 63870
rect 59166 63858 59218 63870
rect 61182 63858 61234 63870
rect 68350 63858 68402 63870
rect 71374 63858 71426 63870
rect 71934 63922 71986 63934
rect 71934 63858 71986 63870
rect 72606 63922 72658 63934
rect 72606 63858 72658 63870
rect 75070 63922 75122 63934
rect 75070 63858 75122 63870
rect 77086 63922 77138 63934
rect 77086 63858 77138 63870
rect 77982 63922 78034 63934
rect 77982 63858 78034 63870
rect 78990 63922 79042 63934
rect 81790 63922 81842 63934
rect 81554 63870 81566 63922
rect 81618 63870 81630 63922
rect 78990 63858 79042 63870
rect 81790 63858 81842 63870
rect 82126 63922 82178 63934
rect 82126 63858 82178 63870
rect 83246 63922 83298 63934
rect 83918 63922 83970 63934
rect 83458 63870 83470 63922
rect 83522 63870 83534 63922
rect 83246 63858 83298 63870
rect 83918 63858 83970 63870
rect 85150 63922 85202 63934
rect 85150 63858 85202 63870
rect 86046 63922 86098 63934
rect 86046 63858 86098 63870
rect 86270 63922 86322 63934
rect 86270 63858 86322 63870
rect 86606 63922 86658 63934
rect 86606 63858 86658 63870
rect 89294 63922 89346 63934
rect 90750 63922 90802 63934
rect 92990 63922 93042 63934
rect 89618 63870 89630 63922
rect 89682 63870 89694 63922
rect 90066 63870 90078 63922
rect 90130 63870 90142 63922
rect 91298 63870 91310 63922
rect 91362 63870 91374 63922
rect 92306 63870 92318 63922
rect 92370 63870 92382 63922
rect 94322 63870 94334 63922
rect 94386 63870 94398 63922
rect 96002 63870 96014 63922
rect 96066 63870 96078 63922
rect 89294 63858 89346 63870
rect 90750 63858 90802 63870
rect 92990 63858 93042 63870
rect 53454 63810 53506 63822
rect 52434 63758 52446 63810
rect 52498 63758 52510 63810
rect 53454 63746 53506 63758
rect 84366 63810 84418 63822
rect 84366 63746 84418 63758
rect 86494 63810 86546 63822
rect 86494 63746 86546 63758
rect 87950 63810 88002 63822
rect 87950 63746 88002 63758
rect 95230 63698 95282 63710
rect 95230 63634 95282 63646
rect 95566 63698 95618 63710
rect 95566 63634 95618 63646
rect 1344 63530 98560 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 96638 63530
rect 96690 63478 96742 63530
rect 96794 63478 96846 63530
rect 96898 63478 98560 63530
rect 1344 63444 98560 63478
rect 72046 63362 72098 63374
rect 72046 63298 72098 63310
rect 52670 63250 52722 63262
rect 50082 63198 50094 63250
rect 50146 63198 50158 63250
rect 52210 63198 52222 63250
rect 52274 63198 52286 63250
rect 52670 63186 52722 63198
rect 57486 63250 57538 63262
rect 66222 63250 66274 63262
rect 58258 63198 58270 63250
rect 58322 63198 58334 63250
rect 59490 63198 59502 63250
rect 59554 63198 59566 63250
rect 57486 63186 57538 63198
rect 66222 63186 66274 63198
rect 68126 63250 68178 63262
rect 68126 63186 68178 63198
rect 77310 63250 77362 63262
rect 77310 63186 77362 63198
rect 79326 63250 79378 63262
rect 79326 63186 79378 63198
rect 86158 63250 86210 63262
rect 86158 63186 86210 63198
rect 92206 63250 92258 63262
rect 92206 63186 92258 63198
rect 96126 63250 96178 63262
rect 96126 63186 96178 63198
rect 55358 63138 55410 63150
rect 58382 63138 58434 63150
rect 59614 63138 59666 63150
rect 49410 63086 49422 63138
rect 49474 63086 49486 63138
rect 54114 63086 54126 63138
rect 54178 63086 54190 63138
rect 54450 63086 54462 63138
rect 54514 63086 54526 63138
rect 55682 63086 55694 63138
rect 55746 63086 55758 63138
rect 56690 63086 56702 63138
rect 56754 63086 56766 63138
rect 58146 63086 58158 63138
rect 58210 63086 58222 63138
rect 59378 63086 59390 63138
rect 59442 63086 59454 63138
rect 55358 63074 55410 63086
rect 58382 63074 58434 63086
rect 59614 63074 59666 63086
rect 62414 63138 62466 63150
rect 62414 63074 62466 63086
rect 67902 63138 67954 63150
rect 67902 63074 67954 63086
rect 68238 63138 68290 63150
rect 68238 63074 68290 63086
rect 68462 63138 68514 63150
rect 68462 63074 68514 63086
rect 70142 63138 70194 63150
rect 70142 63074 70194 63086
rect 71486 63138 71538 63150
rect 71486 63074 71538 63086
rect 71934 63138 71986 63150
rect 71934 63074 71986 63086
rect 72158 63138 72210 63150
rect 76414 63138 76466 63150
rect 81006 63138 81058 63150
rect 83022 63138 83074 63150
rect 72706 63086 72718 63138
rect 72770 63086 72782 63138
rect 77746 63086 77758 63138
rect 77810 63086 77822 63138
rect 78530 63086 78542 63138
rect 78594 63086 78606 63138
rect 79650 63086 79662 63138
rect 79714 63086 79726 63138
rect 80098 63086 80110 63138
rect 80162 63086 80174 63138
rect 81554 63086 81566 63138
rect 81618 63086 81630 63138
rect 82338 63086 82350 63138
rect 82402 63086 82414 63138
rect 72158 63074 72210 63086
rect 76414 63074 76466 63086
rect 81006 63074 81058 63086
rect 83022 63074 83074 63086
rect 84254 63138 84306 63150
rect 84254 63074 84306 63086
rect 86270 63138 86322 63150
rect 89518 63138 89570 63150
rect 86482 63086 86494 63138
rect 86546 63086 86558 63138
rect 88386 63086 88398 63138
rect 88450 63086 88462 63138
rect 88834 63086 88846 63138
rect 88898 63086 88910 63138
rect 90066 63086 90078 63138
rect 90130 63086 90142 63138
rect 91186 63086 91198 63138
rect 91250 63086 91262 63138
rect 86270 63074 86322 63086
rect 89518 63074 89570 63086
rect 1822 63026 1874 63038
rect 1822 62962 1874 62974
rect 53678 63026 53730 63038
rect 58830 63026 58882 63038
rect 54674 62974 54686 63026
rect 54738 62974 54750 63026
rect 53678 62962 53730 62974
rect 58830 62962 58882 62974
rect 60062 63026 60114 63038
rect 60062 62962 60114 62974
rect 61966 63026 62018 63038
rect 61966 62962 62018 62974
rect 62302 63026 62354 63038
rect 69246 63026 69298 63038
rect 67442 62974 67454 63026
rect 67506 62974 67518 63026
rect 62302 62962 62354 62974
rect 69246 62962 69298 62974
rect 73838 63026 73890 63038
rect 73838 62962 73890 62974
rect 75854 63026 75906 63038
rect 83582 63026 83634 63038
rect 78754 62974 78766 63026
rect 78818 62974 78830 63026
rect 75854 62962 75906 62974
rect 83582 62962 83634 62974
rect 83806 63026 83858 63038
rect 83806 62962 83858 62974
rect 85822 63026 85874 63038
rect 85822 62962 85874 62974
rect 86046 63026 86098 63038
rect 86046 62962 86098 62974
rect 88062 63026 88114 63038
rect 88062 62962 88114 62974
rect 94334 63026 94386 63038
rect 94334 62962 94386 62974
rect 95006 63026 95058 63038
rect 95006 62962 95058 62974
rect 95118 63026 95170 63038
rect 95118 62962 95170 62974
rect 2158 62914 2210 62926
rect 2158 62850 2210 62862
rect 58606 62914 58658 62926
rect 58606 62850 58658 62862
rect 59838 62914 59890 62926
rect 59838 62850 59890 62862
rect 62190 62914 62242 62926
rect 62190 62850 62242 62862
rect 62974 62914 63026 62926
rect 62974 62850 63026 62862
rect 63422 62914 63474 62926
rect 63422 62850 63474 62862
rect 65886 62914 65938 62926
rect 65886 62850 65938 62862
rect 67118 62914 67170 62926
rect 67118 62850 67170 62862
rect 69806 62914 69858 62926
rect 69806 62850 69858 62862
rect 70702 62914 70754 62926
rect 70702 62850 70754 62862
rect 71710 62914 71762 62926
rect 83918 62914 83970 62926
rect 76402 62862 76414 62914
rect 76466 62862 76478 62914
rect 80322 62862 80334 62914
rect 80386 62862 80398 62914
rect 71710 62850 71762 62862
rect 83918 62850 83970 62862
rect 85150 62914 85202 62926
rect 85150 62850 85202 62862
rect 86942 62914 86994 62926
rect 86942 62850 86994 62862
rect 87390 62914 87442 62926
rect 91758 62914 91810 62926
rect 89058 62862 89070 62914
rect 89122 62862 89134 62914
rect 87390 62850 87442 62862
rect 91758 62850 91810 62862
rect 93662 62914 93714 62926
rect 93662 62850 93714 62862
rect 93998 62914 94050 62926
rect 93998 62850 94050 62862
rect 94222 62914 94274 62926
rect 94222 62850 94274 62862
rect 94782 62914 94834 62926
rect 94782 62850 94834 62862
rect 95678 62914 95730 62926
rect 95678 62850 95730 62862
rect 1344 62746 98560 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 81278 62746
rect 81330 62694 81382 62746
rect 81434 62694 81486 62746
rect 81538 62694 98560 62746
rect 1344 62660 98560 62694
rect 56702 62578 56754 62590
rect 56702 62514 56754 62526
rect 57598 62578 57650 62590
rect 57598 62514 57650 62526
rect 59278 62578 59330 62590
rect 59278 62514 59330 62526
rect 59502 62578 59554 62590
rect 59502 62514 59554 62526
rect 60286 62578 60338 62590
rect 60286 62514 60338 62526
rect 61966 62578 62018 62590
rect 61966 62514 62018 62526
rect 63310 62578 63362 62590
rect 63310 62514 63362 62526
rect 63982 62578 64034 62590
rect 78430 62578 78482 62590
rect 75394 62526 75406 62578
rect 75458 62526 75470 62578
rect 63982 62514 64034 62526
rect 78430 62514 78482 62526
rect 81566 62578 81618 62590
rect 81566 62514 81618 62526
rect 82462 62578 82514 62590
rect 82462 62514 82514 62526
rect 84366 62578 84418 62590
rect 84366 62514 84418 62526
rect 86270 62578 86322 62590
rect 86270 62514 86322 62526
rect 86606 62578 86658 62590
rect 86606 62514 86658 62526
rect 87614 62578 87666 62590
rect 90290 62526 90302 62578
rect 90354 62526 90366 62578
rect 87614 62514 87666 62526
rect 1822 62466 1874 62478
rect 1822 62402 1874 62414
rect 48750 62466 48802 62478
rect 57822 62466 57874 62478
rect 52658 62414 52670 62466
rect 52722 62414 52734 62466
rect 48750 62402 48802 62414
rect 57822 62402 57874 62414
rect 62190 62466 62242 62478
rect 62190 62402 62242 62414
rect 62414 62466 62466 62478
rect 62414 62402 62466 62414
rect 62974 62466 63026 62478
rect 62974 62402 63026 62414
rect 63198 62466 63250 62478
rect 63198 62402 63250 62414
rect 74846 62466 74898 62478
rect 79438 62466 79490 62478
rect 77522 62414 77534 62466
rect 77586 62414 77598 62466
rect 74846 62402 74898 62414
rect 79438 62402 79490 62414
rect 79774 62466 79826 62478
rect 79774 62402 79826 62414
rect 81342 62466 81394 62478
rect 81342 62402 81394 62414
rect 81902 62466 81954 62478
rect 81902 62402 81954 62414
rect 82798 62466 82850 62478
rect 82798 62402 82850 62414
rect 84590 62466 84642 62478
rect 84590 62402 84642 62414
rect 85150 62466 85202 62478
rect 85150 62402 85202 62414
rect 87278 62466 87330 62478
rect 87278 62402 87330 62414
rect 87502 62466 87554 62478
rect 87502 62402 87554 62414
rect 87838 62466 87890 62478
rect 87838 62402 87890 62414
rect 89294 62466 89346 62478
rect 89294 62402 89346 62414
rect 90750 62466 90802 62478
rect 90750 62402 90802 62414
rect 48414 62354 48466 62366
rect 55806 62354 55858 62366
rect 55346 62302 55358 62354
rect 55410 62302 55422 62354
rect 48414 62290 48466 62302
rect 55806 62290 55858 62302
rect 57374 62354 57426 62366
rect 57374 62290 57426 62302
rect 57934 62354 57986 62366
rect 57934 62290 57986 62302
rect 58606 62354 58658 62366
rect 58606 62290 58658 62302
rect 59166 62354 59218 62366
rect 59166 62290 59218 62302
rect 61854 62354 61906 62366
rect 61854 62290 61906 62302
rect 63534 62354 63586 62366
rect 72046 62354 72098 62366
rect 75406 62354 75458 62366
rect 78094 62354 78146 62366
rect 66322 62302 66334 62354
rect 66386 62302 66398 62354
rect 69906 62302 69918 62354
rect 69970 62302 69982 62354
rect 70130 62302 70142 62354
rect 70194 62302 70206 62354
rect 71026 62302 71038 62354
rect 71090 62302 71102 62354
rect 72482 62302 72494 62354
rect 72546 62302 72558 62354
rect 75730 62302 75742 62354
rect 75794 62302 75806 62354
rect 63534 62290 63586 62302
rect 72046 62290 72098 62302
rect 75406 62290 75458 62302
rect 78094 62290 78146 62302
rect 81678 62354 81730 62366
rect 81678 62290 81730 62302
rect 83246 62354 83298 62366
rect 83246 62290 83298 62302
rect 83694 62354 83746 62366
rect 83694 62290 83746 62302
rect 84702 62354 84754 62366
rect 86382 62354 86434 62366
rect 86034 62302 86046 62354
rect 86098 62302 86110 62354
rect 84702 62290 84754 62302
rect 86382 62290 86434 62302
rect 86494 62354 86546 62366
rect 89618 62302 89630 62354
rect 89682 62302 89694 62354
rect 90178 62302 90190 62354
rect 90242 62302 90254 62354
rect 91522 62302 91534 62354
rect 91586 62302 91598 62354
rect 92306 62302 92318 62354
rect 92370 62302 92382 62354
rect 93650 62302 93662 62354
rect 93714 62302 93726 62354
rect 86494 62290 86546 62302
rect 47854 62242 47906 62254
rect 47854 62178 47906 62190
rect 59950 62242 60002 62254
rect 59950 62178 60002 62190
rect 65774 62242 65826 62254
rect 71486 62242 71538 62254
rect 67106 62190 67118 62242
rect 67170 62190 67182 62242
rect 69234 62190 69246 62242
rect 69298 62190 69310 62242
rect 65774 62178 65826 62190
rect 71486 62178 71538 62190
rect 78878 62242 78930 62254
rect 78878 62178 78930 62190
rect 80222 62242 80274 62254
rect 80222 62178 80274 62190
rect 88286 62242 88338 62254
rect 88286 62178 88338 62190
rect 93102 62242 93154 62254
rect 94322 62190 94334 62242
rect 94386 62190 94398 62242
rect 96450 62190 96462 62242
rect 96514 62190 96526 62242
rect 93102 62178 93154 62190
rect 1344 61962 98560 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 96638 61962
rect 96690 61910 96742 61962
rect 96794 61910 96846 61962
rect 96898 61910 98560 61962
rect 1344 61876 98560 61910
rect 55134 61794 55186 61806
rect 55134 61730 55186 61742
rect 70590 61794 70642 61806
rect 74162 61742 74174 61794
rect 74226 61742 74238 61794
rect 82674 61742 82686 61794
rect 82738 61791 82750 61794
rect 83122 61791 83134 61794
rect 82738 61745 83134 61791
rect 82738 61742 82750 61745
rect 83122 61742 83134 61745
rect 83186 61742 83198 61794
rect 70590 61730 70642 61742
rect 48862 61682 48914 61694
rect 48862 61618 48914 61630
rect 58606 61682 58658 61694
rect 58606 61618 58658 61630
rect 65998 61682 66050 61694
rect 65998 61618 66050 61630
rect 67902 61682 67954 61694
rect 67902 61618 67954 61630
rect 68462 61682 68514 61694
rect 68462 61618 68514 61630
rect 69246 61682 69298 61694
rect 69246 61618 69298 61630
rect 71598 61682 71650 61694
rect 80446 61682 80498 61694
rect 72482 61630 72494 61682
rect 72546 61630 72558 61682
rect 74274 61630 74286 61682
rect 74338 61630 74350 61682
rect 71598 61618 71650 61630
rect 80446 61618 80498 61630
rect 82238 61682 82290 61694
rect 82238 61618 82290 61630
rect 82686 61682 82738 61694
rect 82686 61618 82738 61630
rect 83806 61682 83858 61694
rect 83806 61618 83858 61630
rect 85710 61682 85762 61694
rect 85710 61618 85762 61630
rect 86270 61682 86322 61694
rect 86270 61618 86322 61630
rect 87614 61682 87666 61694
rect 87614 61618 87666 61630
rect 88846 61682 88898 61694
rect 88846 61618 88898 61630
rect 89182 61682 89234 61694
rect 89182 61618 89234 61630
rect 93214 61682 93266 61694
rect 96786 61630 96798 61682
rect 96850 61630 96862 61682
rect 93214 61618 93266 61630
rect 49758 61570 49810 61582
rect 58942 61570 58994 61582
rect 66558 61570 66610 61582
rect 50418 61518 50430 61570
rect 50482 61518 50494 61570
rect 62290 61518 62302 61570
rect 62354 61518 62366 61570
rect 62738 61518 62750 61570
rect 62802 61518 62814 61570
rect 64082 61518 64094 61570
rect 64146 61518 64158 61570
rect 64866 61518 64878 61570
rect 64930 61518 64942 61570
rect 49758 61506 49810 61518
rect 58942 61506 58994 61518
rect 66558 61506 66610 61518
rect 67454 61570 67506 61582
rect 67454 61506 67506 61518
rect 68126 61570 68178 61582
rect 74398 61570 74450 61582
rect 70242 61518 70254 61570
rect 70306 61518 70318 61570
rect 71138 61518 71150 61570
rect 71202 61518 71214 61570
rect 72258 61518 72270 61570
rect 72322 61518 72334 61570
rect 73938 61518 73950 61570
rect 74002 61518 74014 61570
rect 68126 61506 68178 61518
rect 74398 61506 74450 61518
rect 75182 61570 75234 61582
rect 75182 61506 75234 61518
rect 75406 61570 75458 61582
rect 75406 61506 75458 61518
rect 75630 61570 75682 61582
rect 75630 61506 75682 61518
rect 75854 61570 75906 61582
rect 75854 61506 75906 61518
rect 77310 61570 77362 61582
rect 78990 61570 79042 61582
rect 78530 61518 78542 61570
rect 78594 61518 78606 61570
rect 77310 61506 77362 61518
rect 78990 61506 79042 61518
rect 79886 61570 79938 61582
rect 79886 61506 79938 61518
rect 80670 61570 80722 61582
rect 80670 61506 80722 61518
rect 80782 61570 80834 61582
rect 83470 61570 83522 61582
rect 81666 61518 81678 61570
rect 81730 61518 81742 61570
rect 80782 61506 80834 61518
rect 83470 61506 83522 61518
rect 83694 61570 83746 61582
rect 83694 61506 83746 61518
rect 85262 61570 85314 61582
rect 85262 61506 85314 61518
rect 85486 61570 85538 61582
rect 85486 61506 85538 61518
rect 85934 61570 85986 61582
rect 85934 61506 85986 61518
rect 89630 61570 89682 61582
rect 93874 61518 93886 61570
rect 93938 61518 93950 61570
rect 89630 61506 89682 61518
rect 55022 61458 55074 61470
rect 50306 61406 50318 61458
rect 50370 61406 50382 61458
rect 55022 61394 55074 61406
rect 55694 61458 55746 61470
rect 55694 61394 55746 61406
rect 59166 61458 59218 61470
rect 59166 61394 59218 61406
rect 59278 61458 59330 61470
rect 59278 61394 59330 61406
rect 60174 61458 60226 61470
rect 60174 61394 60226 61406
rect 61854 61458 61906 61470
rect 63310 61458 63362 61470
rect 62850 61406 62862 61458
rect 62914 61406 62926 61458
rect 61854 61394 61906 61406
rect 63310 61394 63362 61406
rect 67678 61458 67730 61470
rect 67678 61394 67730 61406
rect 70030 61458 70082 61470
rect 70030 61394 70082 61406
rect 70478 61458 70530 61470
rect 79550 61458 79602 61470
rect 72818 61406 72830 61458
rect 72882 61406 72894 61458
rect 70478 61394 70530 61406
rect 79550 61394 79602 61406
rect 80334 61458 80386 61470
rect 80334 61394 80386 61406
rect 81454 61458 81506 61470
rect 81454 61394 81506 61406
rect 83918 61458 83970 61470
rect 94658 61406 94670 61458
rect 94722 61406 94734 61458
rect 83918 61394 83970 61406
rect 49422 61346 49474 61358
rect 49422 61282 49474 61294
rect 51102 61346 51154 61358
rect 51102 61282 51154 61294
rect 53342 61346 53394 61358
rect 53342 61282 53394 61294
rect 55134 61346 55186 61358
rect 55134 61282 55186 61294
rect 56142 61346 56194 61358
rect 56142 61282 56194 61294
rect 59726 61346 59778 61358
rect 59726 61282 59778 61294
rect 65550 61346 65602 61358
rect 65550 61282 65602 61294
rect 66894 61346 66946 61358
rect 66894 61282 66946 61294
rect 75966 61346 76018 61358
rect 75966 61282 76018 61294
rect 76302 61346 76354 61358
rect 76302 61282 76354 61294
rect 77870 61346 77922 61358
rect 77870 61282 77922 61294
rect 79662 61346 79714 61358
rect 79662 61282 79714 61294
rect 84366 61346 84418 61358
rect 84366 61282 84418 61294
rect 86718 61346 86770 61358
rect 86718 61282 86770 61294
rect 87166 61346 87218 61358
rect 87166 61282 87218 61294
rect 1344 61178 98560 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 81278 61178
rect 81330 61126 81382 61178
rect 81434 61126 81486 61178
rect 81538 61126 98560 61178
rect 1344 61092 98560 61126
rect 56254 61010 56306 61022
rect 66670 61010 66722 61022
rect 62402 60958 62414 61010
rect 62466 60958 62478 61010
rect 56254 60946 56306 60958
rect 66670 60946 66722 60958
rect 69246 61010 69298 61022
rect 88510 61010 88562 61022
rect 85810 60958 85822 61010
rect 85874 60958 85886 61010
rect 69246 60946 69298 60958
rect 88510 60946 88562 60958
rect 90638 61010 90690 61022
rect 90638 60946 90690 60958
rect 48414 60898 48466 60910
rect 48414 60834 48466 60846
rect 48750 60898 48802 60910
rect 55470 60898 55522 60910
rect 50866 60846 50878 60898
rect 50930 60846 50942 60898
rect 48750 60834 48802 60846
rect 55470 60834 55522 60846
rect 65326 60898 65378 60910
rect 68238 60898 68290 60910
rect 67218 60846 67230 60898
rect 67282 60846 67294 60898
rect 65326 60834 65378 60846
rect 68238 60834 68290 60846
rect 68574 60898 68626 60910
rect 68574 60834 68626 60846
rect 70142 60898 70194 60910
rect 70142 60834 70194 60846
rect 70478 60898 70530 60910
rect 70478 60834 70530 60846
rect 71038 60898 71090 60910
rect 71038 60834 71090 60846
rect 71374 60898 71426 60910
rect 71374 60834 71426 60846
rect 72606 60898 72658 60910
rect 72606 60834 72658 60846
rect 79326 60898 79378 60910
rect 79326 60834 79378 60846
rect 79662 60898 79714 60910
rect 82350 60898 82402 60910
rect 80546 60846 80558 60898
rect 80610 60846 80622 60898
rect 79662 60834 79714 60846
rect 82350 60834 82402 60846
rect 82798 60898 82850 60910
rect 82798 60834 82850 60846
rect 84142 60898 84194 60910
rect 84142 60834 84194 60846
rect 50094 60786 50146 60798
rect 55246 60786 55298 60798
rect 50754 60734 50766 60786
rect 50818 60734 50830 60786
rect 50094 60722 50146 60734
rect 55246 60722 55298 60734
rect 55582 60786 55634 60798
rect 55582 60722 55634 60734
rect 56142 60786 56194 60798
rect 56142 60722 56194 60734
rect 56478 60786 56530 60798
rect 63086 60786 63138 60798
rect 67566 60786 67618 60798
rect 61842 60734 61854 60786
rect 61906 60734 61918 60786
rect 62178 60734 62190 60786
rect 62242 60734 62254 60786
rect 63634 60734 63646 60786
rect 63698 60734 63710 60786
rect 64530 60734 64542 60786
rect 64594 60734 64606 60786
rect 56478 60722 56530 60734
rect 63086 60722 63138 60734
rect 67566 60722 67618 60734
rect 69358 60786 69410 60798
rect 80222 60786 80274 60798
rect 72146 60734 72158 60786
rect 72210 60734 72222 60786
rect 78754 60734 78766 60786
rect 78818 60734 78830 60786
rect 69358 60722 69410 60734
rect 80222 60722 80274 60734
rect 81342 60786 81394 60798
rect 81342 60722 81394 60734
rect 83246 60786 83298 60798
rect 83246 60722 83298 60734
rect 84254 60786 84306 60798
rect 89742 60786 89794 60798
rect 85138 60734 85150 60786
rect 85202 60734 85214 60786
rect 85586 60734 85598 60786
rect 85650 60734 85662 60786
rect 86370 60734 86382 60786
rect 86434 60734 86446 60786
rect 87042 60734 87054 60786
rect 87106 60734 87118 60786
rect 87938 60734 87950 60786
rect 88002 60734 88014 60786
rect 95778 60734 95790 60786
rect 95842 60734 95854 60786
rect 84254 60722 84306 60734
rect 89742 60722 89794 60734
rect 51438 60674 51490 60686
rect 51438 60610 51490 60622
rect 51886 60674 51938 60686
rect 51886 60610 51938 60622
rect 57374 60674 57426 60686
rect 57374 60610 57426 60622
rect 57822 60674 57874 60686
rect 57822 60610 57874 60622
rect 61406 60674 61458 60686
rect 61406 60610 61458 60622
rect 65886 60674 65938 60686
rect 65886 60610 65938 60622
rect 66222 60674 66274 60686
rect 81902 60674 81954 60686
rect 76738 60622 76750 60674
rect 76802 60622 76814 60674
rect 66222 60610 66274 60622
rect 81902 60610 81954 60622
rect 84814 60674 84866 60686
rect 84814 60610 84866 60622
rect 89294 60674 89346 60686
rect 93538 60622 93550 60674
rect 93602 60622 93614 60674
rect 89294 60610 89346 60622
rect 49758 60562 49810 60574
rect 69246 60562 69298 60574
rect 65874 60510 65886 60562
rect 65938 60559 65950 60562
rect 66546 60559 66558 60562
rect 65938 60513 66558 60559
rect 65938 60510 65950 60513
rect 66546 60510 66558 60513
rect 66610 60510 66622 60562
rect 49758 60498 49810 60510
rect 69246 60498 69298 60510
rect 81454 60562 81506 60574
rect 81454 60498 81506 60510
rect 84142 60562 84194 60574
rect 84142 60498 84194 60510
rect 1344 60394 98560 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 96638 60394
rect 96690 60342 96742 60394
rect 96794 60342 96846 60394
rect 96898 60342 98560 60394
rect 1344 60308 98560 60342
rect 57262 60226 57314 60238
rect 72718 60226 72770 60238
rect 66098 60174 66110 60226
rect 66162 60223 66174 60226
rect 66770 60223 66782 60226
rect 66162 60177 66782 60223
rect 66162 60174 66174 60177
rect 66770 60174 66782 60177
rect 66834 60174 66846 60226
rect 57262 60162 57314 60174
rect 72718 60162 72770 60174
rect 72942 60226 72994 60238
rect 74946 60174 74958 60226
rect 75010 60174 75022 60226
rect 72942 60162 72994 60174
rect 67230 60114 67282 60126
rect 49074 60062 49086 60114
rect 49138 60062 49150 60114
rect 51202 60062 51214 60114
rect 51266 60062 51278 60114
rect 56578 60062 56590 60114
rect 56642 60062 56654 60114
rect 67230 60050 67282 60062
rect 68462 60114 68514 60126
rect 75854 60114 75906 60126
rect 71474 60062 71486 60114
rect 71538 60062 71550 60114
rect 68462 60050 68514 60062
rect 75854 60050 75906 60062
rect 83134 60114 83186 60126
rect 83134 60050 83186 60062
rect 83582 60114 83634 60126
rect 83582 60050 83634 60062
rect 84030 60114 84082 60126
rect 84030 60050 84082 60062
rect 89070 60114 89122 60126
rect 96450 60062 96462 60114
rect 96514 60062 96526 60114
rect 89070 60050 89122 60062
rect 51774 60002 51826 60014
rect 48402 59950 48414 60002
rect 48466 59950 48478 60002
rect 51774 59938 51826 59950
rect 52782 60002 52834 60014
rect 64430 60002 64482 60014
rect 67678 60002 67730 60014
rect 53666 59950 53678 60002
rect 53730 59950 53742 60002
rect 62850 59950 62862 60002
rect 62914 59950 62926 60002
rect 63634 59950 63646 60002
rect 63698 59950 63710 60002
rect 65090 59950 65102 60002
rect 65154 59950 65166 60002
rect 65538 59950 65550 60002
rect 65602 59950 65614 60002
rect 52782 59938 52834 59950
rect 64430 59938 64482 59950
rect 67678 59938 67730 59950
rect 68014 60002 68066 60014
rect 68014 59938 68066 59950
rect 69470 60002 69522 60014
rect 69470 59938 69522 59950
rect 71934 60002 71986 60014
rect 80894 60002 80946 60014
rect 92206 60002 92258 60014
rect 72482 59950 72494 60002
rect 72546 59950 72558 60002
rect 73938 59950 73950 60002
rect 74002 59950 74014 60002
rect 74498 59950 74510 60002
rect 74562 59950 74574 60002
rect 75282 59950 75294 60002
rect 75346 59950 75358 60002
rect 79762 59950 79774 60002
rect 79826 59950 79838 60002
rect 80210 59950 80222 60002
rect 80274 59950 80286 60002
rect 81666 59950 81678 60002
rect 81730 59950 81742 60002
rect 82450 59950 82462 60002
rect 82514 59950 82526 60002
rect 85586 59950 85598 60002
rect 85650 59950 85662 60002
rect 86034 59950 86046 60002
rect 86098 59950 86110 60002
rect 87490 59950 87502 60002
rect 87554 59950 87566 60002
rect 88386 59950 88398 60002
rect 88450 59950 88462 60002
rect 71934 59938 71986 59950
rect 80894 59938 80946 59950
rect 92206 59938 92258 59950
rect 92542 60002 92594 60014
rect 97694 60002 97746 60014
rect 93538 59950 93550 60002
rect 93602 59950 93614 60002
rect 94322 59950 94334 60002
rect 94386 59950 94398 60002
rect 92542 59938 92594 59950
rect 97694 59938 97746 59950
rect 57262 59890 57314 59902
rect 54450 59838 54462 59890
rect 54514 59838 54526 59890
rect 57262 59826 57314 59838
rect 57374 59890 57426 59902
rect 57374 59826 57426 59838
rect 58382 59890 58434 59902
rect 58382 59826 58434 59838
rect 58494 59890 58546 59902
rect 65886 59890 65938 59902
rect 64866 59838 64878 59890
rect 64930 59838 64942 59890
rect 58494 59826 58546 59838
rect 65886 59826 65938 59838
rect 66782 59890 66834 59902
rect 66782 59826 66834 59838
rect 69806 59890 69858 59902
rect 69806 59826 69858 59838
rect 70478 59890 70530 59902
rect 70478 59826 70530 59838
rect 70814 59890 70866 59902
rect 70814 59826 70866 59838
rect 73054 59890 73106 59902
rect 76414 59890 76466 59902
rect 78206 59890 78258 59902
rect 74050 59838 74062 59890
rect 74114 59838 74126 59890
rect 77634 59838 77646 59890
rect 77698 59838 77710 59890
rect 73054 59826 73106 59838
rect 76414 59826 76466 59838
rect 78206 59826 78258 59838
rect 78542 59890 78594 59902
rect 78542 59826 78594 59838
rect 79438 59890 79490 59902
rect 84478 59890 84530 59902
rect 80434 59838 80446 59890
rect 80498 59838 80510 59890
rect 79438 59826 79490 59838
rect 84478 59826 84530 59838
rect 85262 59890 85314 59902
rect 86718 59890 86770 59902
rect 86258 59838 86270 59890
rect 86322 59838 86334 59890
rect 85262 59826 85314 59838
rect 86718 59826 86770 59838
rect 97022 59890 97074 59902
rect 97022 59826 97074 59838
rect 97134 59890 97186 59902
rect 97134 59826 97186 59838
rect 97358 59890 97410 59902
rect 97358 59826 97410 59838
rect 98030 59890 98082 59902
rect 98030 59826 98082 59838
rect 58158 59778 58210 59790
rect 58158 59714 58210 59726
rect 58942 59778 58994 59790
rect 58942 59714 58994 59726
rect 61742 59778 61794 59790
rect 61742 59714 61794 59726
rect 62190 59778 62242 59790
rect 62190 59714 62242 59726
rect 66334 59778 66386 59790
rect 66334 59714 66386 59726
rect 67902 59778 67954 59790
rect 67902 59714 67954 59726
rect 77310 59778 77362 59790
rect 77310 59714 77362 59726
rect 89406 59778 89458 59790
rect 89406 59714 89458 59726
rect 89854 59778 89906 59790
rect 89854 59714 89906 59726
rect 92318 59778 92370 59790
rect 92318 59714 92370 59726
rect 97918 59778 97970 59790
rect 97918 59714 97970 59726
rect 1344 59610 98560 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 81278 59610
rect 81330 59558 81382 59610
rect 81434 59558 81486 59610
rect 81538 59558 98560 59610
rect 1344 59524 98560 59558
rect 48750 59442 48802 59454
rect 48750 59378 48802 59390
rect 58158 59442 58210 59454
rect 58158 59378 58210 59390
rect 63870 59442 63922 59454
rect 70590 59442 70642 59454
rect 80334 59442 80386 59454
rect 67890 59390 67902 59442
rect 67954 59390 67966 59442
rect 71138 59390 71150 59442
rect 71202 59390 71214 59442
rect 75506 59390 75518 59442
rect 75570 59390 75582 59442
rect 63870 59378 63922 59390
rect 70590 59378 70642 59390
rect 80334 59378 80386 59390
rect 81230 59442 81282 59454
rect 81230 59378 81282 59390
rect 82126 59442 82178 59454
rect 82126 59378 82178 59390
rect 83134 59442 83186 59454
rect 83134 59378 83186 59390
rect 83470 59442 83522 59454
rect 83470 59378 83522 59390
rect 84366 59442 84418 59454
rect 84366 59378 84418 59390
rect 94222 59442 94274 59454
rect 94222 59378 94274 59390
rect 97134 59442 97186 59454
rect 97134 59378 97186 59390
rect 47854 59330 47906 59342
rect 57598 59330 57650 59342
rect 50306 59278 50318 59330
rect 50370 59278 50382 59330
rect 54562 59278 54574 59330
rect 54626 59278 54638 59330
rect 47854 59266 47906 59278
rect 57598 59266 57650 59278
rect 58382 59330 58434 59342
rect 58382 59266 58434 59278
rect 58494 59330 58546 59342
rect 58494 59266 58546 59278
rect 63086 59330 63138 59342
rect 63086 59266 63138 59278
rect 69358 59330 69410 59342
rect 69358 59266 69410 59278
rect 74398 59330 74450 59342
rect 74398 59266 74450 59278
rect 76974 59330 77026 59342
rect 76974 59266 77026 59278
rect 78094 59330 78146 59342
rect 78094 59266 78146 59278
rect 78990 59330 79042 59342
rect 78990 59266 79042 59278
rect 89630 59330 89682 59342
rect 89630 59266 89682 59278
rect 94446 59330 94498 59342
rect 94446 59266 94498 59278
rect 94558 59330 94610 59342
rect 94558 59266 94610 59278
rect 95566 59330 95618 59342
rect 95566 59266 95618 59278
rect 95790 59330 95842 59342
rect 95790 59266 95842 59278
rect 46958 59218 47010 59230
rect 57710 59218 57762 59230
rect 62862 59218 62914 59230
rect 47618 59166 47630 59218
rect 47682 59166 47694 59218
rect 48514 59166 48526 59218
rect 48578 59166 48590 59218
rect 49522 59166 49534 59218
rect 49586 59166 49598 59218
rect 53778 59166 53790 59218
rect 53842 59166 53854 59218
rect 59602 59166 59614 59218
rect 59666 59166 59678 59218
rect 46958 59154 47010 59166
rect 57710 59154 57762 59166
rect 62862 59154 62914 59166
rect 63198 59218 63250 59230
rect 63198 59154 63250 59166
rect 63646 59218 63698 59230
rect 63646 59154 63698 59166
rect 63982 59218 64034 59230
rect 72046 59218 72098 59230
rect 65874 59166 65886 59218
rect 65938 59166 65950 59218
rect 66882 59166 66894 59218
rect 66946 59166 66958 59218
rect 67330 59166 67342 59218
rect 67394 59166 67406 59218
rect 68114 59166 68126 59218
rect 68178 59166 68190 59218
rect 68562 59166 68574 59218
rect 68626 59166 68638 59218
rect 70354 59166 70366 59218
rect 70418 59166 70430 59218
rect 71362 59166 71374 59218
rect 71426 59166 71438 59218
rect 63982 59154 64034 59166
rect 72046 59154 72098 59166
rect 72606 59218 72658 59230
rect 75854 59218 75906 59230
rect 79326 59218 79378 59230
rect 75506 59166 75518 59218
rect 75570 59166 75582 59218
rect 78418 59166 78430 59218
rect 78482 59166 78494 59218
rect 72606 59154 72658 59166
rect 75854 59154 75906 59166
rect 79326 59154 79378 59166
rect 89518 59218 89570 59230
rect 89518 59154 89570 59166
rect 89854 59218 89906 59230
rect 89854 59154 89906 59166
rect 95902 59218 95954 59230
rect 95902 59154 95954 59166
rect 53006 59106 53058 59118
rect 58942 59106 58994 59118
rect 64542 59106 64594 59118
rect 52434 59054 52446 59106
rect 52498 59054 52510 59106
rect 56690 59054 56702 59106
rect 56754 59054 56766 59106
rect 60274 59054 60286 59106
rect 60338 59054 60350 59106
rect 62402 59054 62414 59106
rect 62466 59054 62478 59106
rect 53006 59042 53058 59054
rect 58942 59042 58994 59054
rect 64542 59042 64594 59054
rect 68910 59106 68962 59118
rect 68910 59042 68962 59054
rect 78206 59106 78258 59118
rect 78206 59042 78258 59054
rect 79774 59106 79826 59118
rect 79774 59042 79826 59054
rect 81678 59106 81730 59118
rect 81678 59042 81730 59054
rect 82574 59106 82626 59118
rect 82574 59042 82626 59054
rect 83918 59106 83970 59118
rect 83918 59042 83970 59054
rect 84814 59106 84866 59118
rect 84814 59042 84866 59054
rect 85262 59106 85314 59118
rect 85262 59042 85314 59054
rect 85710 59106 85762 59118
rect 85710 59042 85762 59054
rect 91758 59106 91810 59118
rect 91758 59042 91810 59054
rect 96350 59106 96402 59118
rect 96350 59042 96402 59054
rect 57598 58994 57650 59006
rect 82450 58942 82462 58994
rect 82514 58991 82526 58994
rect 83906 58991 83918 58994
rect 82514 58945 83918 58991
rect 82514 58942 82526 58945
rect 83906 58942 83918 58945
rect 83970 58942 83982 58994
rect 57598 58930 57650 58942
rect 1344 58826 98560 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 96638 58826
rect 96690 58774 96742 58826
rect 96794 58774 96846 58826
rect 96898 58774 98560 58826
rect 1344 58740 98560 58774
rect 64990 58658 65042 58670
rect 51090 58606 51102 58658
rect 51154 58655 51166 58658
rect 51650 58655 51662 58658
rect 51154 58609 51662 58655
rect 51154 58606 51166 58609
rect 51650 58606 51662 58609
rect 51714 58606 51726 58658
rect 69122 58606 69134 58658
rect 69186 58655 69198 58658
rect 69794 58655 69806 58658
rect 69186 58609 69806 58655
rect 69186 58606 69198 58609
rect 69794 58606 69806 58609
rect 69858 58606 69870 58658
rect 83458 58606 83470 58658
rect 83522 58655 83534 58658
rect 84466 58655 84478 58658
rect 83522 58609 84478 58655
rect 83522 58606 83534 58609
rect 84466 58606 84478 58609
rect 84530 58606 84542 58658
rect 64990 58594 65042 58606
rect 47966 58546 48018 58558
rect 47966 58482 48018 58494
rect 51102 58546 51154 58558
rect 51102 58482 51154 58494
rect 51998 58546 52050 58558
rect 69358 58546 69410 58558
rect 58034 58494 58046 58546
rect 58098 58494 58110 58546
rect 61394 58494 61406 58546
rect 61458 58494 61470 58546
rect 63522 58494 63534 58546
rect 63586 58494 63598 58546
rect 51998 58482 52050 58494
rect 69358 58482 69410 58494
rect 70254 58546 70306 58558
rect 78878 58546 78930 58558
rect 72258 58494 72270 58546
rect 72322 58494 72334 58546
rect 70254 58482 70306 58494
rect 78878 58482 78930 58494
rect 80222 58546 80274 58558
rect 80222 58482 80274 58494
rect 81118 58546 81170 58558
rect 81118 58482 81170 58494
rect 83134 58546 83186 58558
rect 83134 58482 83186 58494
rect 83582 58546 83634 58558
rect 83582 58482 83634 58494
rect 84142 58546 84194 58558
rect 84142 58482 84194 58494
rect 84478 58546 84530 58558
rect 84478 58482 84530 58494
rect 85150 58546 85202 58558
rect 88498 58494 88510 58546
rect 88562 58494 88574 58546
rect 90626 58494 90638 58546
rect 90690 58494 90702 58546
rect 85150 58482 85202 58494
rect 49422 58434 49474 58446
rect 48514 58382 48526 58434
rect 48578 58382 48590 58434
rect 49422 58370 49474 58382
rect 49758 58434 49810 58446
rect 54350 58434 54402 58446
rect 58494 58434 58546 58446
rect 50530 58382 50542 58434
rect 50594 58382 50606 58434
rect 55234 58382 55246 58434
rect 55298 58382 55310 58434
rect 49758 58370 49810 58382
rect 54350 58370 54402 58382
rect 58494 58370 58546 58382
rect 59838 58434 59890 58446
rect 59838 58370 59890 58382
rect 60286 58434 60338 58446
rect 65102 58434 65154 58446
rect 64194 58382 64206 58434
rect 64258 58382 64270 58434
rect 60286 58370 60338 58382
rect 65102 58370 65154 58382
rect 68238 58434 68290 58446
rect 68238 58370 68290 58382
rect 68574 58434 68626 58446
rect 75630 58434 75682 58446
rect 72146 58382 72158 58434
rect 72210 58382 72222 58434
rect 73490 58382 73502 58434
rect 73554 58382 73566 58434
rect 74050 58382 74062 58434
rect 74114 58382 74126 58434
rect 74610 58382 74622 58434
rect 74674 58382 74686 58434
rect 68574 58370 68626 58382
rect 75630 58370 75682 58382
rect 76078 58434 76130 58446
rect 76078 58370 76130 58382
rect 79774 58434 79826 58446
rect 95678 58434 95730 58446
rect 91410 58382 91422 58434
rect 91474 58382 91486 58434
rect 79774 58370 79826 58382
rect 95678 58370 95730 58382
rect 54462 58322 54514 58334
rect 50418 58270 50430 58322
rect 50482 58270 50494 58322
rect 54462 58258 54514 58270
rect 54686 58322 54738 58334
rect 60622 58322 60674 58334
rect 55906 58270 55918 58322
rect 55970 58270 55982 58322
rect 54686 58258 54738 58270
rect 60622 58258 60674 58270
rect 65550 58322 65602 58334
rect 65550 58258 65602 58270
rect 65774 58322 65826 58334
rect 65774 58258 65826 58270
rect 65886 58322 65938 58334
rect 65886 58258 65938 58270
rect 70814 58322 70866 58334
rect 70814 58258 70866 58270
rect 71150 58322 71202 58334
rect 73278 58322 73330 58334
rect 75406 58322 75458 58334
rect 71810 58270 71822 58322
rect 71874 58270 71886 58322
rect 73602 58270 73614 58322
rect 73666 58270 73678 58322
rect 71150 58258 71202 58270
rect 73278 58258 73330 58270
rect 75406 58258 75458 58270
rect 77310 58322 77362 58334
rect 77310 58258 77362 58270
rect 77646 58322 77698 58334
rect 77646 58258 77698 58270
rect 78206 58322 78258 58334
rect 78206 58258 78258 58270
rect 78318 58322 78370 58334
rect 78318 58258 78370 58270
rect 81566 58322 81618 58334
rect 81566 58258 81618 58270
rect 87726 58322 87778 58334
rect 87726 58258 87778 58270
rect 87838 58322 87890 58334
rect 87838 58258 87890 58270
rect 94894 58322 94946 58334
rect 94894 58258 94946 58270
rect 96462 58322 96514 58334
rect 96462 58258 96514 58270
rect 48750 58210 48802 58222
rect 48750 58146 48802 58158
rect 51662 58210 51714 58222
rect 51662 58146 51714 58158
rect 52670 58210 52722 58222
rect 52670 58146 52722 58158
rect 53454 58210 53506 58222
rect 53454 58146 53506 58158
rect 60510 58210 60562 58222
rect 60510 58146 60562 58158
rect 64990 58210 65042 58222
rect 64990 58146 65042 58158
rect 66446 58210 66498 58222
rect 66446 58146 66498 58158
rect 66894 58210 66946 58222
rect 66894 58146 66946 58158
rect 69806 58210 69858 58222
rect 69806 58146 69858 58158
rect 72830 58210 72882 58222
rect 72830 58146 72882 58158
rect 75294 58210 75346 58222
rect 75294 58146 75346 58158
rect 75854 58210 75906 58222
rect 75854 58146 75906 58158
rect 76526 58210 76578 58222
rect 76526 58146 76578 58158
rect 78542 58210 78594 58222
rect 78542 58146 78594 58158
rect 79326 58210 79378 58222
rect 79326 58146 79378 58158
rect 80670 58210 80722 58222
rect 80670 58146 80722 58158
rect 82126 58210 82178 58222
rect 82126 58146 82178 58158
rect 86830 58210 86882 58222
rect 86830 58146 86882 58158
rect 87278 58210 87330 58222
rect 87278 58146 87330 58158
rect 88062 58210 88114 58222
rect 88062 58146 88114 58158
rect 91982 58210 92034 58222
rect 91982 58146 92034 58158
rect 92430 58210 92482 58222
rect 92430 58146 92482 58158
rect 93214 58210 93266 58222
rect 93214 58146 93266 58158
rect 94558 58210 94610 58222
rect 94558 58146 94610 58158
rect 94782 58210 94834 58222
rect 94782 58146 94834 58158
rect 95342 58210 95394 58222
rect 95342 58146 95394 58158
rect 95566 58210 95618 58222
rect 95566 58146 95618 58158
rect 96126 58210 96178 58222
rect 96126 58146 96178 58158
rect 96350 58210 96402 58222
rect 96350 58146 96402 58158
rect 96910 58210 96962 58222
rect 96910 58146 96962 58158
rect 97358 58210 97410 58222
rect 97358 58146 97410 58158
rect 1344 58042 98560 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 81278 58042
rect 81330 57990 81382 58042
rect 81434 57990 81486 58042
rect 81538 57990 98560 58042
rect 1344 57956 98560 57990
rect 65326 57874 65378 57886
rect 51426 57822 51438 57874
rect 51490 57822 51502 57874
rect 65326 57810 65378 57822
rect 65550 57874 65602 57886
rect 65550 57810 65602 57822
rect 66110 57874 66162 57886
rect 66110 57810 66162 57822
rect 69582 57874 69634 57886
rect 69582 57810 69634 57822
rect 70030 57874 70082 57886
rect 70030 57810 70082 57822
rect 70366 57874 70418 57886
rect 70366 57810 70418 57822
rect 73502 57874 73554 57886
rect 77422 57874 77474 57886
rect 76178 57822 76190 57874
rect 76242 57822 76254 57874
rect 73502 57810 73554 57822
rect 77422 57810 77474 57822
rect 78878 57874 78930 57886
rect 78878 57810 78930 57822
rect 82014 57874 82066 57886
rect 82014 57810 82066 57822
rect 97582 57874 97634 57886
rect 97582 57810 97634 57822
rect 53118 57762 53170 57774
rect 50642 57710 50654 57762
rect 50706 57710 50718 57762
rect 53118 57698 53170 57710
rect 57598 57762 57650 57774
rect 57598 57698 57650 57710
rect 57710 57762 57762 57774
rect 65662 57762 65714 57774
rect 60946 57710 60958 57762
rect 61010 57710 61022 57762
rect 57710 57698 57762 57710
rect 65662 57698 65714 57710
rect 73614 57762 73666 57774
rect 73614 57698 73666 57710
rect 74846 57762 74898 57774
rect 76862 57762 76914 57774
rect 75842 57710 75854 57762
rect 75906 57710 75918 57762
rect 74846 57698 74898 57710
rect 76862 57698 76914 57710
rect 76974 57762 77026 57774
rect 76974 57698 77026 57710
rect 78542 57762 78594 57774
rect 78542 57698 78594 57710
rect 79438 57762 79490 57774
rect 79438 57698 79490 57710
rect 79550 57762 79602 57774
rect 79550 57698 79602 57710
rect 80334 57762 80386 57774
rect 80334 57698 80386 57710
rect 80446 57762 80498 57774
rect 80446 57698 80498 57710
rect 80670 57762 80722 57774
rect 80670 57698 80722 57710
rect 81342 57762 81394 57774
rect 81342 57698 81394 57710
rect 81454 57762 81506 57774
rect 88286 57762 88338 57774
rect 84690 57710 84702 57762
rect 84754 57710 84766 57762
rect 81454 57698 81506 57710
rect 88286 57698 88338 57710
rect 88398 57762 88450 57774
rect 88398 57698 88450 57710
rect 92766 57762 92818 57774
rect 92766 57698 92818 57710
rect 92878 57762 92930 57774
rect 97246 57762 97298 57774
rect 94322 57710 94334 57762
rect 94386 57710 94398 57762
rect 92878 57698 92930 57710
rect 97246 57698 97298 57710
rect 97358 57762 97410 57774
rect 97358 57698 97410 57710
rect 51774 57650 51826 57662
rect 50754 57598 50766 57650
rect 50818 57598 50830 57650
rect 51774 57586 51826 57598
rect 53006 57650 53058 57662
rect 53006 57586 53058 57598
rect 53342 57650 53394 57662
rect 67006 57650 67058 57662
rect 53778 57598 53790 57650
rect 53842 57598 53854 57650
rect 60386 57598 60398 57650
rect 60450 57598 60462 57650
rect 53342 57586 53394 57598
rect 67006 57586 67058 57598
rect 67566 57650 67618 57662
rect 67566 57586 67618 57598
rect 71598 57650 71650 57662
rect 71598 57586 71650 57598
rect 71822 57650 71874 57662
rect 71822 57586 71874 57598
rect 74286 57650 74338 57662
rect 74286 57586 74338 57598
rect 74734 57650 74786 57662
rect 74734 57586 74786 57598
rect 75070 57650 75122 57662
rect 82910 57650 82962 57662
rect 88622 57650 88674 57662
rect 93102 57650 93154 57662
rect 75730 57598 75742 57650
rect 75794 57598 75806 57650
rect 84018 57598 84030 57650
rect 84082 57598 84094 57650
rect 84466 57598 84478 57650
rect 84530 57598 84542 57650
rect 85250 57598 85262 57650
rect 85314 57598 85326 57650
rect 85922 57598 85934 57650
rect 85986 57598 85998 57650
rect 86818 57598 86830 57650
rect 86882 57598 86894 57650
rect 91410 57598 91422 57650
rect 91474 57598 91486 57650
rect 92194 57598 92206 57650
rect 92258 57598 92270 57650
rect 93650 57598 93662 57650
rect 93714 57598 93726 57650
rect 75070 57586 75122 57598
rect 82910 57586 82962 57598
rect 88622 57586 88674 57598
rect 93102 57586 93154 57598
rect 52222 57538 52274 57550
rect 64766 57538 64818 57550
rect 54562 57486 54574 57538
rect 54626 57486 54638 57538
rect 56690 57486 56702 57538
rect 56754 57486 56766 57538
rect 52222 57474 52274 57486
rect 64766 57474 64818 57486
rect 68014 57538 68066 57550
rect 68014 57474 68066 57486
rect 68798 57538 68850 57550
rect 68798 57474 68850 57486
rect 70814 57538 70866 57550
rect 70814 57474 70866 57486
rect 72606 57538 72658 57550
rect 72606 57474 72658 57486
rect 77870 57538 77922 57550
rect 77870 57474 77922 57486
rect 82574 57538 82626 57550
rect 82574 57474 82626 57486
rect 83694 57538 83746 57550
rect 83694 57474 83746 57486
rect 87502 57538 87554 57550
rect 97918 57538 97970 57550
rect 89282 57486 89294 57538
rect 89346 57486 89358 57538
rect 96450 57486 96462 57538
rect 96514 57486 96526 57538
rect 87502 57474 87554 57486
rect 97918 57474 97970 57486
rect 49646 57426 49698 57438
rect 49646 57362 49698 57374
rect 49982 57426 50034 57438
rect 49982 57362 50034 57374
rect 57598 57426 57650 57438
rect 73502 57426 73554 57438
rect 72146 57374 72158 57426
rect 72210 57374 72222 57426
rect 57598 57362 57650 57374
rect 73502 57362 73554 57374
rect 74062 57426 74114 57438
rect 74062 57362 74114 57374
rect 79550 57426 79602 57438
rect 79550 57362 79602 57374
rect 81454 57426 81506 57438
rect 81454 57362 81506 57374
rect 1344 57258 98560 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 96638 57258
rect 96690 57206 96742 57258
rect 96794 57206 96846 57258
rect 96898 57206 98560 57258
rect 1344 57172 98560 57206
rect 57374 57090 57426 57102
rect 57374 57026 57426 57038
rect 88622 57090 88674 57102
rect 88622 57026 88674 57038
rect 70142 56978 70194 56990
rect 49074 56926 49086 56978
rect 49138 56926 49150 56978
rect 51202 56926 51214 56978
rect 51266 56926 51278 56978
rect 54338 56926 54350 56978
rect 54402 56926 54414 56978
rect 56466 56926 56478 56978
rect 56530 56926 56542 56978
rect 62178 56926 62190 56978
rect 62242 56926 62254 56978
rect 64306 56926 64318 56978
rect 64370 56926 64382 56978
rect 70142 56914 70194 56926
rect 70590 56978 70642 56990
rect 70590 56914 70642 56926
rect 72718 56978 72770 56990
rect 73614 56978 73666 56990
rect 73042 56926 73054 56978
rect 73106 56926 73118 56978
rect 72718 56914 72770 56926
rect 73614 56914 73666 56926
rect 76414 56978 76466 56990
rect 87390 56978 87442 56990
rect 78978 56926 78990 56978
rect 79042 56926 79054 56978
rect 81106 56926 81118 56978
rect 81170 56926 81182 56978
rect 76414 56914 76466 56926
rect 87390 56914 87442 56926
rect 87950 56978 88002 56990
rect 92194 56926 92206 56978
rect 92258 56926 92270 56978
rect 94994 56926 95006 56978
rect 95058 56926 95070 56978
rect 97122 56926 97134 56978
rect 97186 56926 97198 56978
rect 87950 56914 88002 56926
rect 57486 56866 57538 56878
rect 48402 56814 48414 56866
rect 48466 56814 48478 56866
rect 53554 56814 53566 56866
rect 53618 56814 53630 56866
rect 57486 56802 57538 56814
rect 57934 56866 57986 56878
rect 68574 56866 68626 56878
rect 61506 56814 61518 56866
rect 61570 56814 61582 56866
rect 68114 56814 68126 56866
rect 68178 56814 68190 56866
rect 57934 56802 57986 56814
rect 68574 56802 68626 56814
rect 69694 56866 69746 56878
rect 73838 56866 73890 56878
rect 81566 56866 81618 56878
rect 84030 56866 84082 56878
rect 71810 56814 71822 56866
rect 71874 56814 71886 56866
rect 74162 56814 74174 56866
rect 74226 56814 74238 56866
rect 78194 56814 78206 56866
rect 78258 56814 78270 56866
rect 83234 56814 83246 56866
rect 83298 56814 83310 56866
rect 69694 56802 69746 56814
rect 73838 56802 73890 56814
rect 81566 56802 81618 56814
rect 84030 56802 84082 56814
rect 88510 56866 88562 56878
rect 93438 56866 93490 56878
rect 89394 56814 89406 56866
rect 89458 56814 89470 56866
rect 94322 56814 94334 56866
rect 94386 56814 94398 56866
rect 88510 56802 88562 56814
rect 93438 56802 93490 56814
rect 57374 56754 57426 56766
rect 57374 56690 57426 56702
rect 58270 56754 58322 56766
rect 58270 56690 58322 56702
rect 74958 56754 75010 56766
rect 74958 56690 75010 56702
rect 75294 56754 75346 56766
rect 75294 56690 75346 56702
rect 75966 56754 76018 56766
rect 75966 56690 76018 56702
rect 81790 56754 81842 56766
rect 81790 56690 81842 56702
rect 81902 56754 81954 56766
rect 88622 56754 88674 56766
rect 83458 56702 83470 56754
rect 83522 56702 83534 56754
rect 90066 56702 90078 56754
rect 90130 56702 90142 56754
rect 81902 56690 81954 56702
rect 88622 56690 88674 56702
rect 51662 56642 51714 56654
rect 51662 56578 51714 56590
rect 52670 56642 52722 56654
rect 52670 56578 52722 56590
rect 58158 56642 58210 56654
rect 58158 56578 58210 56590
rect 58718 56642 58770 56654
rect 58718 56578 58770 56590
rect 59166 56642 59218 56654
rect 59166 56578 59218 56590
rect 64766 56642 64818 56654
rect 64766 56578 64818 56590
rect 65214 56642 65266 56654
rect 65214 56578 65266 56590
rect 69358 56642 69410 56654
rect 69358 56578 69410 56590
rect 71150 56642 71202 56654
rect 75854 56642 75906 56654
rect 71586 56590 71598 56642
rect 71650 56590 71662 56642
rect 71150 56578 71202 56590
rect 75854 56578 75906 56590
rect 77198 56642 77250 56654
rect 77198 56578 77250 56590
rect 77646 56642 77698 56654
rect 77646 56578 77698 56590
rect 82574 56642 82626 56654
rect 82574 56578 82626 56590
rect 84366 56642 84418 56654
rect 84366 56578 84418 56590
rect 85150 56642 85202 56654
rect 85150 56578 85202 56590
rect 93102 56642 93154 56654
rect 93102 56578 93154 56590
rect 93326 56642 93378 56654
rect 93326 56578 93378 56590
rect 97582 56642 97634 56654
rect 97582 56578 97634 56590
rect 1344 56474 98560 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 81278 56474
rect 81330 56422 81382 56474
rect 81434 56422 81486 56474
rect 81538 56422 98560 56474
rect 1344 56388 98560 56422
rect 50654 56306 50706 56318
rect 50654 56242 50706 56254
rect 57374 56306 57426 56318
rect 57374 56242 57426 56254
rect 68014 56306 68066 56318
rect 68014 56242 68066 56254
rect 68238 56306 68290 56318
rect 68238 56242 68290 56254
rect 70926 56306 70978 56318
rect 70926 56242 70978 56254
rect 71486 56306 71538 56318
rect 71486 56242 71538 56254
rect 71934 56306 71986 56318
rect 71934 56242 71986 56254
rect 72494 56306 72546 56318
rect 72494 56242 72546 56254
rect 73726 56306 73778 56318
rect 73726 56242 73778 56254
rect 73950 56306 74002 56318
rect 73950 56242 74002 56254
rect 75406 56306 75458 56318
rect 75406 56242 75458 56254
rect 77310 56306 77362 56318
rect 77310 56242 77362 56254
rect 77870 56306 77922 56318
rect 77870 56242 77922 56254
rect 79438 56306 79490 56318
rect 79438 56242 79490 56254
rect 80334 56306 80386 56318
rect 80334 56242 80386 56254
rect 88622 56306 88674 56318
rect 88622 56242 88674 56254
rect 90526 56306 90578 56318
rect 90526 56242 90578 56254
rect 57598 56194 57650 56206
rect 51426 56142 51438 56194
rect 51490 56142 51502 56194
rect 57598 56130 57650 56142
rect 57710 56194 57762 56206
rect 57710 56130 57762 56142
rect 60846 56194 60898 56206
rect 60846 56130 60898 56142
rect 60958 56194 61010 56206
rect 60958 56130 61010 56142
rect 65550 56194 65602 56206
rect 65550 56130 65602 56142
rect 67454 56194 67506 56206
rect 67454 56130 67506 56142
rect 67566 56194 67618 56206
rect 67566 56130 67618 56142
rect 72382 56194 72434 56206
rect 72382 56130 72434 56142
rect 73502 56194 73554 56206
rect 73502 56130 73554 56142
rect 74510 56194 74562 56206
rect 74510 56130 74562 56142
rect 74846 56194 74898 56206
rect 74846 56130 74898 56142
rect 76302 56194 76354 56206
rect 76302 56130 76354 56142
rect 76638 56194 76690 56206
rect 76638 56130 76690 56142
rect 77422 56194 77474 56206
rect 77422 56130 77474 56142
rect 78878 56194 78930 56206
rect 78878 56130 78930 56142
rect 79998 56194 80050 56206
rect 79998 56130 80050 56142
rect 88286 56194 88338 56206
rect 88286 56130 88338 56142
rect 88398 56194 88450 56206
rect 88398 56130 88450 56142
rect 89630 56194 89682 56206
rect 89630 56130 89682 56142
rect 89742 56194 89794 56206
rect 89742 56130 89794 56142
rect 90302 56194 90354 56206
rect 90302 56130 90354 56142
rect 65326 56082 65378 56094
rect 56466 56030 56478 56082
rect 56530 56030 56542 56082
rect 61618 56030 61630 56082
rect 61682 56030 61694 56082
rect 65326 56018 65378 56030
rect 65662 56082 65714 56094
rect 65662 56018 65714 56030
rect 66110 56082 66162 56094
rect 66110 56018 66162 56030
rect 68350 56082 68402 56094
rect 68350 56018 68402 56030
rect 68910 56082 68962 56094
rect 68910 56018 68962 56030
rect 75742 56082 75794 56094
rect 75742 56018 75794 56030
rect 77086 56082 77138 56094
rect 77086 56018 77138 56030
rect 78766 56082 78818 56094
rect 87502 56082 87554 56094
rect 82786 56030 82798 56082
rect 82850 56030 82862 56082
rect 78766 56018 78818 56030
rect 87502 56018 87554 56030
rect 90638 56082 90690 56094
rect 92306 56030 92318 56082
rect 92370 56030 92382 56082
rect 90638 56018 90690 56030
rect 58158 55970 58210 55982
rect 97246 55970 97298 55982
rect 62402 55918 62414 55970
rect 62466 55918 62478 55970
rect 64530 55918 64542 55970
rect 64594 55918 64606 55970
rect 84018 55918 84030 55970
rect 84082 55918 84094 55970
rect 96226 55918 96238 55970
rect 96290 55918 96302 55970
rect 58158 55906 58210 55918
rect 97246 55906 97298 55918
rect 60958 55858 61010 55870
rect 60958 55794 61010 55806
rect 67454 55858 67506 55870
rect 67454 55794 67506 55806
rect 72494 55858 72546 55870
rect 72494 55794 72546 55806
rect 74062 55858 74114 55870
rect 74062 55794 74114 55806
rect 78878 55858 78930 55870
rect 78878 55794 78930 55806
rect 89742 55858 89794 55870
rect 89742 55794 89794 55806
rect 1344 55690 98560 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 96638 55690
rect 96690 55638 96742 55690
rect 96794 55638 96846 55690
rect 96898 55638 98560 55690
rect 1344 55604 98560 55638
rect 78990 55522 79042 55534
rect 78990 55458 79042 55470
rect 92318 55410 92370 55422
rect 96910 55410 96962 55422
rect 51202 55358 51214 55410
rect 51266 55358 51278 55410
rect 54450 55358 54462 55410
rect 54514 55358 54526 55410
rect 56578 55358 56590 55410
rect 56642 55358 56654 55410
rect 80546 55358 80558 55410
rect 80610 55358 80622 55410
rect 82674 55358 82686 55410
rect 82738 55358 82750 55410
rect 88162 55358 88174 55410
rect 88226 55358 88238 55410
rect 89730 55358 89742 55410
rect 89794 55358 89806 55410
rect 91858 55358 91870 55410
rect 91922 55358 91934 55410
rect 94322 55358 94334 55410
rect 94386 55358 94398 55410
rect 96450 55358 96462 55410
rect 96514 55358 96526 55410
rect 92318 55346 92370 55358
rect 96910 55346 96962 55358
rect 60622 55298 60674 55310
rect 77758 55298 77810 55310
rect 48402 55246 48414 55298
rect 48466 55246 48478 55298
rect 53778 55246 53790 55298
rect 53842 55246 53854 55298
rect 68562 55246 68574 55298
rect 68626 55246 68638 55298
rect 70690 55246 70702 55298
rect 70754 55246 70766 55298
rect 72034 55246 72046 55298
rect 72098 55246 72110 55298
rect 72706 55246 72718 55298
rect 72770 55246 72782 55298
rect 74946 55246 74958 55298
rect 75010 55246 75022 55298
rect 60622 55234 60674 55246
rect 77758 55234 77810 55246
rect 78318 55298 78370 55310
rect 79762 55246 79774 55298
rect 79826 55246 79838 55298
rect 83346 55246 83358 55298
rect 83410 55246 83422 55298
rect 84354 55246 84366 55298
rect 84418 55246 84430 55298
rect 85250 55246 85262 55298
rect 85314 55246 85326 55298
rect 89058 55246 89070 55298
rect 89122 55246 89134 55298
rect 93538 55246 93550 55298
rect 93602 55246 93614 55298
rect 78318 55234 78370 55246
rect 51774 55186 51826 55198
rect 49074 55134 49086 55186
rect 49138 55134 49150 55186
rect 51774 55122 51826 55134
rect 52110 55186 52162 55198
rect 52110 55122 52162 55134
rect 52558 55186 52610 55198
rect 52558 55122 52610 55134
rect 61294 55186 61346 55198
rect 61294 55122 61346 55134
rect 62414 55186 62466 55198
rect 73390 55186 73442 55198
rect 77198 55186 77250 55198
rect 63858 55134 63870 55186
rect 63922 55134 63934 55186
rect 76514 55134 76526 55186
rect 76578 55134 76590 55186
rect 62414 55122 62466 55134
rect 73390 55122 73442 55134
rect 77198 55122 77250 55134
rect 78990 55186 79042 55198
rect 83582 55186 83634 55198
rect 78990 55122 79042 55134
rect 79102 55130 79154 55142
rect 57038 55074 57090 55086
rect 57038 55010 57090 55022
rect 62078 55074 62130 55086
rect 62078 55010 62130 55022
rect 62302 55074 62354 55086
rect 70926 55074 70978 55086
rect 68562 55022 68574 55074
rect 68626 55071 68638 55074
rect 68786 55071 68798 55074
rect 68626 55025 68798 55071
rect 68626 55022 68638 55025
rect 68786 55022 68798 55025
rect 68850 55022 68862 55074
rect 62302 55010 62354 55022
rect 70926 55010 70978 55022
rect 71822 55074 71874 55086
rect 86034 55134 86046 55186
rect 86098 55134 86110 55186
rect 83582 55122 83634 55134
rect 75506 55022 75518 55074
rect 75570 55022 75582 55074
rect 79102 55066 79154 55078
rect 84142 55074 84194 55086
rect 71822 55010 71874 55022
rect 84142 55010 84194 55022
rect 1344 54906 98560 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 81278 54906
rect 81330 54854 81382 54906
rect 81434 54854 81486 54906
rect 81538 54854 98560 54906
rect 1344 54820 98560 54854
rect 48750 54738 48802 54750
rect 48750 54674 48802 54686
rect 54350 54738 54402 54750
rect 54350 54674 54402 54686
rect 55470 54738 55522 54750
rect 55470 54674 55522 54686
rect 56702 54738 56754 54750
rect 56702 54674 56754 54686
rect 59726 54738 59778 54750
rect 59726 54674 59778 54686
rect 63982 54738 64034 54750
rect 63982 54674 64034 54686
rect 72270 54738 72322 54750
rect 72270 54674 72322 54686
rect 72606 54738 72658 54750
rect 72606 54674 72658 54686
rect 74958 54738 75010 54750
rect 74958 54674 75010 54686
rect 85598 54738 85650 54750
rect 85598 54674 85650 54686
rect 86046 54738 86098 54750
rect 86046 54674 86098 54686
rect 87502 54738 87554 54750
rect 87502 54674 87554 54686
rect 88510 54738 88562 54750
rect 88510 54674 88562 54686
rect 89294 54738 89346 54750
rect 89294 54674 89346 54686
rect 90862 54738 90914 54750
rect 90862 54674 90914 54686
rect 93102 54738 93154 54750
rect 93102 54674 93154 54686
rect 93886 54738 93938 54750
rect 93886 54674 93938 54686
rect 94670 54738 94722 54750
rect 94670 54674 94722 54686
rect 48414 54626 48466 54638
rect 55694 54626 55746 54638
rect 50866 54574 50878 54626
rect 50930 54574 50942 54626
rect 52882 54574 52894 54626
rect 52946 54574 52958 54626
rect 48414 54562 48466 54574
rect 55694 54562 55746 54574
rect 56478 54626 56530 54638
rect 56478 54562 56530 54574
rect 59950 54626 60002 54638
rect 64206 54626 64258 54638
rect 61394 54574 61406 54626
rect 61458 54574 61470 54626
rect 59950 54562 60002 54574
rect 64206 54562 64258 54574
rect 64318 54626 64370 54638
rect 69134 54626 69186 54638
rect 66434 54574 66446 54626
rect 66498 54574 66510 54626
rect 64318 54562 64370 54574
rect 69134 54562 69186 54574
rect 69470 54626 69522 54638
rect 69470 54562 69522 54574
rect 69918 54626 69970 54638
rect 69918 54562 69970 54574
rect 71150 54626 71202 54638
rect 71150 54562 71202 54574
rect 76414 54626 76466 54638
rect 76414 54562 76466 54574
rect 76750 54626 76802 54638
rect 85262 54626 85314 54638
rect 78418 54574 78430 54626
rect 78482 54574 78494 54626
rect 82562 54574 82574 54626
rect 82626 54574 82638 54626
rect 76750 54562 76802 54574
rect 85262 54562 85314 54574
rect 88286 54626 88338 54638
rect 88286 54562 88338 54574
rect 89518 54626 89570 54638
rect 89518 54562 89570 54574
rect 90302 54626 90354 54638
rect 90302 54562 90354 54574
rect 91086 54626 91138 54638
rect 91086 54562 91138 54574
rect 92766 54626 92818 54638
rect 92766 54562 92818 54574
rect 92878 54626 92930 54638
rect 92878 54562 92930 54574
rect 93550 54626 93602 54638
rect 93550 54562 93602 54574
rect 93662 54626 93714 54638
rect 93662 54562 93714 54574
rect 94446 54626 94498 54638
rect 94446 54562 94498 54574
rect 50206 54514 50258 54526
rect 52110 54514 52162 54526
rect 55022 54514 55074 54526
rect 50978 54462 50990 54514
rect 51042 54462 51054 54514
rect 52770 54462 52782 54514
rect 52834 54462 52846 54514
rect 50206 54450 50258 54462
rect 52110 54450 52162 54462
rect 55022 54450 55074 54462
rect 55806 54514 55858 54526
rect 55806 54450 55858 54462
rect 56366 54514 56418 54526
rect 56366 54450 56418 54462
rect 60062 54514 60114 54526
rect 73838 54514 73890 54526
rect 60722 54462 60734 54514
rect 60786 54462 60798 54514
rect 65650 54462 65662 54514
rect 65714 54462 65726 54514
rect 60062 54450 60114 54462
rect 73838 54450 73890 54462
rect 74062 54514 74114 54526
rect 86830 54514 86882 54526
rect 77746 54462 77758 54514
rect 77810 54462 77822 54514
rect 81778 54462 81790 54514
rect 81842 54462 81854 54514
rect 74062 54450 74114 54462
rect 86830 54450 86882 54462
rect 87390 54514 87442 54526
rect 87390 54450 87442 54462
rect 88174 54514 88226 54526
rect 88174 54450 88226 54462
rect 89630 54514 89682 54526
rect 89630 54450 89682 54462
rect 90078 54514 90130 54526
rect 90078 54450 90130 54462
rect 90414 54514 90466 54526
rect 90414 54450 90466 54462
rect 91198 54514 91250 54526
rect 91198 54450 91250 54462
rect 94334 54514 94386 54526
rect 94334 54450 94386 54462
rect 53454 54402 53506 54414
rect 53454 54338 53506 54350
rect 53902 54402 53954 54414
rect 53902 54338 53954 54350
rect 57374 54402 57426 54414
rect 57374 54338 57426 54350
rect 57822 54402 57874 54414
rect 57822 54338 57874 54350
rect 59278 54402 59330 54414
rect 71710 54402 71762 54414
rect 63522 54350 63534 54402
rect 63586 54350 63598 54402
rect 68562 54350 68574 54402
rect 68626 54350 68638 54402
rect 59278 54338 59330 54350
rect 71710 54338 71762 54350
rect 73390 54402 73442 54414
rect 81342 54402 81394 54414
rect 91646 54402 91698 54414
rect 75394 54350 75406 54402
rect 75458 54350 75470 54402
rect 80546 54350 80558 54402
rect 80610 54350 80622 54402
rect 84690 54350 84702 54402
rect 84754 54350 84766 54402
rect 73390 54338 73442 54350
rect 81342 54338 81394 54350
rect 91646 54338 91698 54350
rect 92094 54402 92146 54414
rect 92094 54338 92146 54350
rect 95006 54402 95058 54414
rect 95006 54338 95058 54350
rect 98030 54402 98082 54414
rect 98030 54338 98082 54350
rect 49870 54290 49922 54302
rect 49870 54226 49922 54238
rect 51774 54290 51826 54302
rect 51774 54226 51826 54238
rect 73614 54290 73666 54302
rect 73614 54226 73666 54238
rect 74510 54290 74562 54302
rect 74510 54226 74562 54238
rect 87502 54290 87554 54302
rect 87502 54226 87554 54238
rect 1344 54122 98560 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 96638 54122
rect 96690 54070 96742 54122
rect 96794 54070 96846 54122
rect 96898 54070 98560 54122
rect 1344 54036 98560 54070
rect 83806 53954 83858 53966
rect 60050 53902 60062 53954
rect 60114 53951 60126 53954
rect 60274 53951 60286 53954
rect 60114 53905 60286 53951
rect 60114 53902 60126 53905
rect 60274 53902 60286 53905
rect 60338 53902 60350 53954
rect 72594 53902 72606 53954
rect 72658 53951 72670 53954
rect 73602 53951 73614 53954
rect 72658 53905 73614 53951
rect 72658 53902 72670 53905
rect 73602 53902 73614 53905
rect 73666 53902 73678 53954
rect 83806 53890 83858 53902
rect 84142 53954 84194 53966
rect 84142 53890 84194 53902
rect 74734 53842 74786 53854
rect 51650 53790 51662 53842
rect 51714 53790 51726 53842
rect 64306 53790 64318 53842
rect 64370 53790 64382 53842
rect 74734 53778 74786 53790
rect 75854 53842 75906 53854
rect 91646 53842 91698 53854
rect 80210 53790 80222 53842
rect 80274 53790 80286 53842
rect 87826 53790 87838 53842
rect 87890 53790 87902 53842
rect 75854 53778 75906 53790
rect 91646 53778 91698 53790
rect 93102 53842 93154 53854
rect 93102 53778 93154 53790
rect 93662 53842 93714 53854
rect 93662 53778 93714 53790
rect 94110 53842 94162 53854
rect 94770 53790 94782 53842
rect 94834 53790 94846 53842
rect 94110 53778 94162 53790
rect 52110 53730 52162 53742
rect 47954 53678 47966 53730
rect 48018 53678 48030 53730
rect 48850 53678 48862 53730
rect 48914 53678 48926 53730
rect 52110 53666 52162 53678
rect 56366 53730 56418 53742
rect 56366 53666 56418 53678
rect 56702 53730 56754 53742
rect 56702 53666 56754 53678
rect 57486 53730 57538 53742
rect 64766 53730 64818 53742
rect 61506 53678 61518 53730
rect 61570 53678 61582 53730
rect 62178 53678 62190 53730
rect 62242 53678 62254 53730
rect 57486 53666 57538 53678
rect 64766 53666 64818 53678
rect 65326 53730 65378 53742
rect 65326 53666 65378 53678
rect 67006 53730 67058 53742
rect 67006 53666 67058 53678
rect 67454 53730 67506 53742
rect 67454 53666 67506 53678
rect 67790 53730 67842 53742
rect 67790 53666 67842 53678
rect 76302 53730 76354 53742
rect 87278 53730 87330 53742
rect 91198 53730 91250 53742
rect 77410 53678 77422 53730
rect 77474 53678 77486 53730
rect 83234 53678 83246 53730
rect 83298 53678 83310 53730
rect 90738 53678 90750 53730
rect 90802 53678 90814 53730
rect 76302 53666 76354 53678
rect 87278 53666 87330 53678
rect 91198 53666 91250 53678
rect 92318 53730 92370 53742
rect 97682 53678 97694 53730
rect 97746 53678 97758 53730
rect 92318 53666 92370 53678
rect 48190 53618 48242 53630
rect 65550 53618 65602 53630
rect 49522 53566 49534 53618
rect 49586 53566 49598 53618
rect 48190 53554 48242 53566
rect 65550 53554 65602 53566
rect 65662 53618 65714 53630
rect 65662 53554 65714 53566
rect 66110 53618 66162 53630
rect 66110 53554 66162 53566
rect 68574 53618 68626 53630
rect 68574 53554 68626 53566
rect 69582 53618 69634 53630
rect 69582 53554 69634 53566
rect 70366 53618 70418 53630
rect 70366 53554 70418 53566
rect 76414 53618 76466 53630
rect 76414 53554 76466 53566
rect 76638 53618 76690 53630
rect 85150 53618 85202 53630
rect 78082 53566 78094 53618
rect 78146 53566 78158 53618
rect 83010 53566 83022 53618
rect 83074 53566 83086 53618
rect 76638 53554 76690 53566
rect 85150 53554 85202 53566
rect 86382 53618 86434 53630
rect 86382 53554 86434 53566
rect 86942 53618 86994 53630
rect 89954 53566 89966 53618
rect 90018 53566 90030 53618
rect 96898 53566 96910 53618
rect 96962 53566 96974 53618
rect 86942 53554 86994 53566
rect 52558 53506 52610 53518
rect 52558 53442 52610 53454
rect 56478 53506 56530 53518
rect 56478 53442 56530 53454
rect 57150 53506 57202 53518
rect 57150 53442 57202 53454
rect 60286 53506 60338 53518
rect 60286 53442 60338 53454
rect 67678 53506 67730 53518
rect 67678 53442 67730 53454
rect 68238 53506 68290 53518
rect 68238 53442 68290 53454
rect 68462 53506 68514 53518
rect 68462 53442 68514 53454
rect 69246 53506 69298 53518
rect 69246 53442 69298 53454
rect 69470 53506 69522 53518
rect 69470 53442 69522 53454
rect 70030 53506 70082 53518
rect 70030 53442 70082 53454
rect 70254 53506 70306 53518
rect 70254 53442 70306 53454
rect 70814 53506 70866 53518
rect 70814 53442 70866 53454
rect 71262 53506 71314 53518
rect 71262 53442 71314 53454
rect 72494 53506 72546 53518
rect 72494 53442 72546 53454
rect 73054 53506 73106 53518
rect 73054 53442 73106 53454
rect 73502 53506 73554 53518
rect 73502 53442 73554 53454
rect 80670 53506 80722 53518
rect 80670 53442 80722 53454
rect 82350 53506 82402 53518
rect 82350 53442 82402 53454
rect 87054 53506 87106 53518
rect 87054 53442 87106 53454
rect 1344 53338 98560 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 81278 53338
rect 81330 53286 81382 53338
rect 81434 53286 81486 53338
rect 81538 53286 98560 53338
rect 1344 53252 98560 53286
rect 52894 53170 52946 53182
rect 52894 53106 52946 53118
rect 61630 53170 61682 53182
rect 61630 53106 61682 53118
rect 61854 53170 61906 53182
rect 61854 53106 61906 53118
rect 62862 53170 62914 53182
rect 62862 53106 62914 53118
rect 63198 53170 63250 53182
rect 63198 53106 63250 53118
rect 63422 53170 63474 53182
rect 63422 53106 63474 53118
rect 65326 53170 65378 53182
rect 65326 53106 65378 53118
rect 65774 53170 65826 53182
rect 65774 53106 65826 53118
rect 70366 53170 70418 53182
rect 70366 53106 70418 53118
rect 71150 53170 71202 53182
rect 71150 53106 71202 53118
rect 72270 53170 72322 53182
rect 72270 53106 72322 53118
rect 75294 53170 75346 53182
rect 75294 53106 75346 53118
rect 75742 53170 75794 53182
rect 75742 53106 75794 53118
rect 77646 53170 77698 53182
rect 77646 53106 77698 53118
rect 78430 53170 78482 53182
rect 78430 53106 78482 53118
rect 78654 53170 78706 53182
rect 78654 53106 78706 53118
rect 79550 53170 79602 53182
rect 79550 53106 79602 53118
rect 83022 53170 83074 53182
rect 83022 53106 83074 53118
rect 89406 53170 89458 53182
rect 89406 53106 89458 53118
rect 89630 53170 89682 53182
rect 89630 53106 89682 53118
rect 90526 53170 90578 53182
rect 90526 53106 90578 53118
rect 92206 53170 92258 53182
rect 92206 53106 92258 53118
rect 95678 53170 95730 53182
rect 95678 53106 95730 53118
rect 98030 53170 98082 53182
rect 98030 53106 98082 53118
rect 62638 53058 62690 53070
rect 62638 52994 62690 53006
rect 63534 53058 63586 53070
rect 63534 52994 63586 53006
rect 64542 53058 64594 53070
rect 89294 53058 89346 53070
rect 67330 53006 67342 53058
rect 67394 53006 67406 53058
rect 70802 53006 70814 53058
rect 70866 53006 70878 53058
rect 87378 53006 87390 53058
rect 87442 53006 87454 53058
rect 64542 52994 64594 53006
rect 89294 52994 89346 53006
rect 94670 53058 94722 53070
rect 94670 52994 94722 53006
rect 95454 53058 95506 53070
rect 95454 52994 95506 53006
rect 96238 53058 96290 53070
rect 96238 52994 96290 53006
rect 61966 52946 62018 52958
rect 49522 52894 49534 52946
rect 49586 52894 49598 52946
rect 61966 52882 62018 52894
rect 62526 52946 62578 52958
rect 73390 52946 73442 52958
rect 66546 52894 66558 52946
rect 66610 52894 66622 52946
rect 62526 52882 62578 52894
rect 73390 52882 73442 52894
rect 78318 52946 78370 52958
rect 78318 52882 78370 52894
rect 79102 52946 79154 52958
rect 90078 52946 90130 52958
rect 88162 52894 88174 52946
rect 88226 52894 88238 52946
rect 79102 52882 79154 52894
rect 90078 52882 90130 52894
rect 94558 52946 94610 52958
rect 94558 52882 94610 52894
rect 95342 52946 95394 52958
rect 95342 52882 95394 52894
rect 96126 52946 96178 52958
rect 96126 52882 96178 52894
rect 96462 52946 96514 52958
rect 96462 52882 96514 52894
rect 97582 52946 97634 52958
rect 97582 52882 97634 52894
rect 61182 52834 61234 52846
rect 50306 52782 50318 52834
rect 50370 52782 50382 52834
rect 52434 52782 52446 52834
rect 52498 52782 52510 52834
rect 61182 52770 61234 52782
rect 63982 52834 64034 52846
rect 71710 52834 71762 52846
rect 74398 52834 74450 52846
rect 90862 52834 90914 52846
rect 69458 52782 69470 52834
rect 69522 52782 69534 52834
rect 73826 52782 73838 52834
rect 73890 52782 73902 52834
rect 85250 52782 85262 52834
rect 85314 52782 85326 52834
rect 63982 52770 64034 52782
rect 71710 52770 71762 52782
rect 74398 52770 74450 52782
rect 90862 52770 90914 52782
rect 92654 52834 92706 52846
rect 92654 52770 92706 52782
rect 93214 52834 93266 52846
rect 93214 52770 93266 52782
rect 93550 52834 93602 52846
rect 93550 52770 93602 52782
rect 93998 52834 94050 52846
rect 93998 52770 94050 52782
rect 97134 52834 97186 52846
rect 97134 52770 97186 52782
rect 94670 52722 94722 52734
rect 94670 52658 94722 52670
rect 1344 52554 98560 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 96638 52554
rect 96690 52502 96742 52554
rect 96794 52502 96846 52554
rect 96898 52502 98560 52554
rect 1344 52468 98560 52502
rect 62178 52334 62190 52386
rect 62242 52383 62254 52386
rect 62626 52383 62638 52386
rect 62242 52337 62638 52383
rect 62242 52334 62254 52337
rect 62626 52334 62638 52337
rect 62690 52334 62702 52386
rect 53342 52274 53394 52286
rect 53342 52210 53394 52222
rect 62190 52274 62242 52286
rect 62190 52210 62242 52222
rect 66334 52274 66386 52286
rect 66334 52210 66386 52222
rect 69806 52274 69858 52286
rect 69806 52210 69858 52222
rect 73502 52274 73554 52286
rect 73502 52210 73554 52222
rect 73950 52274 74002 52286
rect 73950 52210 74002 52222
rect 77646 52274 77698 52286
rect 77646 52210 77698 52222
rect 78766 52274 78818 52286
rect 78766 52210 78818 52222
rect 86046 52274 86098 52286
rect 94770 52222 94782 52274
rect 94834 52222 94846 52274
rect 86046 52210 86098 52222
rect 53790 52162 53842 52174
rect 53790 52098 53842 52110
rect 54574 52162 54626 52174
rect 56254 52162 56306 52174
rect 58718 52162 58770 52174
rect 55010 52110 55022 52162
rect 55074 52110 55086 52162
rect 55346 52110 55358 52162
rect 55410 52110 55422 52162
rect 56578 52110 56590 52162
rect 56642 52110 56654 52162
rect 57586 52110 57598 52162
rect 57650 52110 57662 52162
rect 54574 52098 54626 52110
rect 56254 52098 56306 52110
rect 58718 52098 58770 52110
rect 62638 52162 62690 52174
rect 62638 52098 62690 52110
rect 67006 52162 67058 52174
rect 67006 52098 67058 52110
rect 68126 52162 68178 52174
rect 71262 52162 71314 52174
rect 74734 52162 74786 52174
rect 70130 52110 70142 52162
rect 70194 52110 70206 52162
rect 70690 52110 70702 52162
rect 70754 52110 70766 52162
rect 72034 52110 72046 52162
rect 72098 52110 72110 52162
rect 72818 52110 72830 52162
rect 72882 52110 72894 52162
rect 68126 52098 68178 52110
rect 71262 52098 71314 52110
rect 74734 52098 74786 52110
rect 75742 52162 75794 52174
rect 75742 52098 75794 52110
rect 76302 52162 76354 52174
rect 76302 52098 76354 52110
rect 85486 52162 85538 52174
rect 87502 52162 87554 52174
rect 92430 52162 92482 52174
rect 86370 52110 86382 52162
rect 86434 52110 86446 52162
rect 86930 52110 86942 52162
rect 86994 52110 87006 52162
rect 88274 52110 88286 52162
rect 88338 52110 88350 52162
rect 89170 52110 89182 52162
rect 89234 52110 89246 52162
rect 91186 52110 91198 52162
rect 91250 52110 91262 52162
rect 85486 52098 85538 52110
rect 87502 52098 87554 52110
rect 92430 52098 92482 52110
rect 94334 52162 94386 52174
rect 97682 52110 97694 52162
rect 97746 52110 97758 52162
rect 94334 52098 94386 52110
rect 49310 52050 49362 52062
rect 49310 51986 49362 51998
rect 49646 52050 49698 52062
rect 67118 52050 67170 52062
rect 55570 51998 55582 52050
rect 55634 51998 55646 52050
rect 49646 51986 49698 51998
rect 67118 51986 67170 51998
rect 67790 52050 67842 52062
rect 67790 51986 67842 51998
rect 67902 52050 67954 52062
rect 67902 51986 67954 51998
rect 68462 52050 68514 52062
rect 89854 52050 89906 52062
rect 70802 51998 70814 52050
rect 70866 51998 70878 52050
rect 87042 51998 87054 52050
rect 87106 51998 87118 52050
rect 68462 51986 68514 51998
rect 89854 51986 89906 51998
rect 93326 52050 93378 52062
rect 93326 51986 93378 51998
rect 93438 52050 93490 52062
rect 93438 51986 93490 51998
rect 93998 52050 94050 52062
rect 93998 51986 94050 51998
rect 94110 52050 94162 52062
rect 96898 51998 96910 52050
rect 96962 51998 96974 52050
rect 94110 51986 94162 51998
rect 58270 51938 58322 51950
rect 58270 51874 58322 51886
rect 67342 51938 67394 51950
rect 67342 51874 67394 51886
rect 75070 51938 75122 51950
rect 75070 51874 75122 51886
rect 77198 51938 77250 51950
rect 77198 51874 77250 51886
rect 90190 51938 90242 51950
rect 90190 51874 90242 51886
rect 91422 51938 91474 51950
rect 91422 51874 91474 51886
rect 91870 51938 91922 51950
rect 91870 51874 91922 51886
rect 93102 51938 93154 51950
rect 93102 51874 93154 51886
rect 1344 51770 98560 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 81278 51770
rect 81330 51718 81382 51770
rect 81434 51718 81486 51770
rect 81538 51718 98560 51770
rect 1344 51684 98560 51718
rect 53118 51602 53170 51614
rect 53118 51538 53170 51550
rect 54350 51602 54402 51614
rect 54350 51538 54402 51550
rect 57374 51602 57426 51614
rect 61630 51602 61682 51614
rect 60162 51550 60174 51602
rect 60226 51550 60238 51602
rect 57374 51538 57426 51550
rect 61630 51538 61682 51550
rect 62078 51602 62130 51614
rect 62078 51538 62130 51550
rect 63982 51602 64034 51614
rect 63982 51538 64034 51550
rect 65326 51602 65378 51614
rect 65326 51538 65378 51550
rect 74062 51602 74114 51614
rect 74062 51538 74114 51550
rect 74510 51602 74562 51614
rect 74510 51538 74562 51550
rect 75518 51602 75570 51614
rect 75518 51538 75570 51550
rect 76862 51602 76914 51614
rect 76862 51538 76914 51550
rect 77422 51602 77474 51614
rect 77422 51538 77474 51550
rect 82462 51602 82514 51614
rect 82462 51538 82514 51550
rect 89630 51602 89682 51614
rect 89630 51538 89682 51550
rect 97134 51602 97186 51614
rect 97134 51538 97186 51550
rect 97358 51602 97410 51614
rect 97358 51538 97410 51550
rect 97918 51602 97970 51614
rect 97918 51538 97970 51550
rect 59726 51490 59778 51502
rect 73502 51490 73554 51502
rect 78318 51490 78370 51502
rect 68002 51438 68014 51490
rect 68066 51438 68078 51490
rect 75842 51438 75854 51490
rect 75906 51438 75918 51490
rect 59726 51426 59778 51438
rect 73502 51426 73554 51438
rect 78318 51426 78370 51438
rect 79102 51490 79154 51502
rect 79102 51426 79154 51438
rect 79214 51490 79266 51502
rect 79214 51426 79266 51438
rect 79438 51490 79490 51502
rect 79438 51426 79490 51438
rect 79998 51490 80050 51502
rect 79998 51426 80050 51438
rect 81230 51490 81282 51502
rect 81230 51426 81282 51438
rect 81454 51490 81506 51502
rect 97470 51490 97522 51502
rect 96226 51438 96238 51490
rect 96290 51438 96302 51490
rect 81454 51426 81506 51438
rect 97470 51426 97522 51438
rect 64094 51378 64146 51390
rect 73278 51378 73330 51390
rect 58034 51326 58046 51378
rect 58098 51326 58110 51378
rect 59154 51326 59166 51378
rect 59218 51326 59230 51378
rect 60274 51326 60286 51378
rect 60338 51326 60350 51378
rect 60834 51326 60846 51378
rect 60898 51326 60910 51378
rect 67330 51326 67342 51378
rect 67394 51326 67406 51378
rect 64094 51314 64146 51326
rect 73278 51314 73330 51326
rect 73614 51378 73666 51390
rect 73614 51314 73666 51326
rect 76750 51378 76802 51390
rect 76750 51314 76802 51326
rect 77086 51378 77138 51390
rect 77086 51314 77138 51326
rect 78206 51378 78258 51390
rect 78206 51314 78258 51326
rect 79886 51378 79938 51390
rect 79886 51314 79938 51326
rect 81566 51378 81618 51390
rect 91970 51326 91982 51378
rect 92034 51326 92046 51378
rect 81566 51314 81618 51326
rect 54798 51266 54850 51278
rect 54798 51202 54850 51214
rect 55246 51266 55298 51278
rect 55246 51202 55298 51214
rect 55694 51266 55746 51278
rect 55694 51202 55746 51214
rect 56030 51266 56082 51278
rect 56030 51202 56082 51214
rect 61182 51266 61234 51278
rect 61182 51202 61234 51214
rect 62638 51266 62690 51278
rect 62638 51202 62690 51214
rect 62974 51266 63026 51278
rect 62974 51202 63026 51214
rect 64542 51266 64594 51278
rect 70702 51266 70754 51278
rect 70130 51214 70142 51266
rect 70194 51214 70206 51266
rect 64542 51202 64594 51214
rect 70702 51202 70754 51214
rect 71038 51266 71090 51278
rect 71038 51202 71090 51214
rect 71710 51266 71762 51278
rect 71710 51202 71762 51214
rect 75070 51266 75122 51278
rect 75070 51202 75122 51214
rect 80558 51266 80610 51278
rect 80558 51202 80610 51214
rect 82014 51266 82066 51278
rect 82014 51202 82066 51214
rect 85710 51266 85762 51278
rect 85710 51202 85762 51214
rect 89966 51266 90018 51278
rect 89966 51202 90018 51214
rect 90414 51266 90466 51278
rect 90414 51202 90466 51214
rect 63982 51154 64034 51166
rect 54226 51102 54238 51154
rect 54290 51151 54302 51154
rect 55234 51151 55246 51154
rect 54290 51105 55246 51151
rect 54290 51102 54302 51105
rect 55234 51102 55246 51105
rect 55298 51102 55310 51154
rect 63982 51090 64034 51102
rect 78318 51154 78370 51166
rect 78318 51090 78370 51102
rect 79998 51154 80050 51166
rect 89506 51102 89518 51154
rect 89570 51151 89582 51154
rect 90402 51151 90414 51154
rect 89570 51105 90414 51151
rect 89570 51102 89582 51105
rect 90402 51102 90414 51105
rect 90466 51102 90478 51154
rect 79998 51090 80050 51102
rect 1344 50986 98560 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 96638 50986
rect 96690 50934 96742 50986
rect 96794 50934 96846 50986
rect 96898 50934 98560 50986
rect 1344 50900 98560 50934
rect 93326 50818 93378 50830
rect 65986 50766 65998 50818
rect 66050 50815 66062 50818
rect 66546 50815 66558 50818
rect 66050 50769 66558 50815
rect 66050 50766 66062 50769
rect 66546 50766 66558 50769
rect 66610 50766 66622 50818
rect 93326 50754 93378 50766
rect 58382 50706 58434 50718
rect 58382 50642 58434 50654
rect 58942 50706 58994 50718
rect 58942 50642 58994 50654
rect 59390 50706 59442 50718
rect 59390 50642 59442 50654
rect 59726 50706 59778 50718
rect 59726 50642 59778 50654
rect 60174 50706 60226 50718
rect 65998 50706 66050 50718
rect 64754 50654 64766 50706
rect 64818 50654 64830 50706
rect 60174 50642 60226 50654
rect 65998 50642 66050 50654
rect 69246 50706 69298 50718
rect 73938 50654 73950 50706
rect 74002 50654 74014 50706
rect 80658 50654 80670 50706
rect 80722 50654 80734 50706
rect 97794 50654 97806 50706
rect 97858 50654 97870 50706
rect 69246 50642 69298 50654
rect 51550 50594 51602 50606
rect 51550 50530 51602 50542
rect 53678 50594 53730 50606
rect 56926 50594 56978 50606
rect 75854 50594 75906 50606
rect 83806 50594 83858 50606
rect 55234 50542 55246 50594
rect 55298 50542 55310 50594
rect 56354 50542 56366 50594
rect 56418 50542 56430 50594
rect 57474 50542 57486 50594
rect 57538 50542 57550 50594
rect 58034 50542 58046 50594
rect 58098 50542 58110 50594
rect 61842 50542 61854 50594
rect 61906 50542 61918 50594
rect 71138 50542 71150 50594
rect 71202 50542 71214 50594
rect 74946 50542 74958 50594
rect 75010 50542 75022 50594
rect 79538 50542 79550 50594
rect 79602 50542 79614 50594
rect 53678 50530 53730 50542
rect 56926 50530 56978 50542
rect 75854 50530 75906 50542
rect 83806 50530 83858 50542
rect 91086 50594 91138 50606
rect 91086 50530 91138 50542
rect 92430 50594 92482 50606
rect 92430 50530 92482 50542
rect 93214 50594 93266 50606
rect 93214 50530 93266 50542
rect 93998 50594 94050 50606
rect 94994 50542 95006 50594
rect 95058 50542 95070 50594
rect 93998 50530 94050 50542
rect 50990 50482 51042 50494
rect 50990 50418 51042 50430
rect 52334 50482 52386 50494
rect 52334 50418 52386 50430
rect 52670 50482 52722 50494
rect 52670 50418 52722 50430
rect 54238 50482 54290 50494
rect 65326 50482 65378 50494
rect 62626 50430 62638 50482
rect 62690 50430 62702 50482
rect 54238 50418 54290 50430
rect 65326 50418 65378 50430
rect 70030 50482 70082 50494
rect 77198 50482 77250 50494
rect 71810 50430 71822 50482
rect 71874 50430 71886 50482
rect 70030 50418 70082 50430
rect 77198 50418 77250 50430
rect 85262 50482 85314 50494
rect 85262 50418 85314 50430
rect 85822 50482 85874 50494
rect 85822 50418 85874 50430
rect 87278 50482 87330 50494
rect 87278 50418 87330 50430
rect 88958 50482 89010 50494
rect 88958 50418 89010 50430
rect 89294 50482 89346 50494
rect 89294 50418 89346 50430
rect 89966 50482 90018 50494
rect 89966 50418 90018 50430
rect 90078 50482 90130 50494
rect 90078 50418 90130 50430
rect 91534 50482 91586 50494
rect 91534 50418 91586 50430
rect 91870 50482 91922 50494
rect 91870 50418 91922 50430
rect 94110 50482 94162 50494
rect 95666 50430 95678 50482
rect 95730 50430 95742 50482
rect 94110 50418 94162 50430
rect 51886 50370 51938 50382
rect 51886 50306 51938 50318
rect 52558 50370 52610 50382
rect 52558 50306 52610 50318
rect 53342 50370 53394 50382
rect 53342 50306 53394 50318
rect 53566 50370 53618 50382
rect 53566 50306 53618 50318
rect 54350 50370 54402 50382
rect 54350 50306 54402 50318
rect 54574 50370 54626 50382
rect 65438 50370 65490 50382
rect 57362 50318 57374 50370
rect 57426 50318 57438 50370
rect 54574 50306 54626 50318
rect 65438 50306 65490 50318
rect 65662 50370 65714 50382
rect 65662 50306 65714 50318
rect 66446 50370 66498 50382
rect 66446 50306 66498 50318
rect 69694 50370 69746 50382
rect 69694 50306 69746 50318
rect 69918 50370 69970 50382
rect 69918 50306 69970 50318
rect 70478 50370 70530 50382
rect 70478 50306 70530 50318
rect 75182 50370 75234 50382
rect 75182 50306 75234 50318
rect 76190 50370 76242 50382
rect 76190 50306 76242 50318
rect 89742 50370 89794 50382
rect 89742 50306 89794 50318
rect 90750 50370 90802 50382
rect 90750 50306 90802 50318
rect 90974 50370 91026 50382
rect 90974 50306 91026 50318
rect 91758 50370 91810 50382
rect 91758 50306 91810 50318
rect 93326 50370 93378 50382
rect 93326 50306 93378 50318
rect 94334 50370 94386 50382
rect 94334 50306 94386 50318
rect 1344 50202 98560 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 81278 50202
rect 81330 50150 81382 50202
rect 81434 50150 81486 50202
rect 81538 50150 98560 50202
rect 1344 50116 98560 50150
rect 56702 50034 56754 50046
rect 56702 49970 56754 49982
rect 57598 50034 57650 50046
rect 57598 49970 57650 49982
rect 68350 50034 68402 50046
rect 68350 49970 68402 49982
rect 71934 50034 71986 50046
rect 71934 49970 71986 49982
rect 72158 50034 72210 50046
rect 72158 49970 72210 49982
rect 76414 50034 76466 50046
rect 76414 49970 76466 49982
rect 76862 50034 76914 50046
rect 85038 50034 85090 50046
rect 82338 49982 82350 50034
rect 82402 49982 82414 50034
rect 76862 49970 76914 49982
rect 85038 49970 85090 49982
rect 89406 50034 89458 50046
rect 89406 49970 89458 49982
rect 90190 50034 90242 50046
rect 90190 49970 90242 49982
rect 95566 50034 95618 50046
rect 95566 49970 95618 49982
rect 96126 50034 96178 50046
rect 96126 49970 96178 49982
rect 96350 50034 96402 50046
rect 96350 49970 96402 49982
rect 55582 49922 55634 49934
rect 55582 49858 55634 49870
rect 65550 49922 65602 49934
rect 65550 49858 65602 49870
rect 65662 49922 65714 49934
rect 65662 49858 65714 49870
rect 66334 49922 66386 49934
rect 66334 49858 66386 49870
rect 66894 49922 66946 49934
rect 66894 49858 66946 49870
rect 68910 49922 68962 49934
rect 68910 49858 68962 49870
rect 69358 49922 69410 49934
rect 69358 49858 69410 49870
rect 70590 49922 70642 49934
rect 70590 49858 70642 49870
rect 71486 49922 71538 49934
rect 71486 49858 71538 49870
rect 72270 49922 72322 49934
rect 72270 49858 72322 49870
rect 73390 49922 73442 49934
rect 73390 49858 73442 49870
rect 73726 49922 73778 49934
rect 73726 49858 73778 49870
rect 74286 49922 74338 49934
rect 74286 49858 74338 49870
rect 74622 49922 74674 49934
rect 74622 49858 74674 49870
rect 75182 49922 75234 49934
rect 75182 49858 75234 49870
rect 75518 49922 75570 49934
rect 75518 49858 75570 49870
rect 76078 49922 76130 49934
rect 86494 49922 86546 49934
rect 78306 49870 78318 49922
rect 78370 49870 78382 49922
rect 76078 49858 76130 49870
rect 86494 49858 86546 49870
rect 87614 49922 87666 49934
rect 87614 49858 87666 49870
rect 88398 49922 88450 49934
rect 88398 49858 88450 49870
rect 90302 49922 90354 49934
rect 94782 49922 94834 49934
rect 93314 49870 93326 49922
rect 93378 49870 93390 49922
rect 90302 49858 90354 49870
rect 94782 49858 94834 49870
rect 94894 49922 94946 49934
rect 94894 49858 94946 49870
rect 95454 49922 95506 49934
rect 95454 49858 95506 49870
rect 95790 49922 95842 49934
rect 95790 49858 95842 49870
rect 96462 49922 96514 49934
rect 96462 49858 96514 49870
rect 97358 49922 97410 49934
rect 97358 49858 97410 49870
rect 97470 49922 97522 49934
rect 97470 49858 97522 49870
rect 57486 49810 57538 49822
rect 51874 49758 51886 49810
rect 51938 49758 51950 49810
rect 55346 49758 55358 49810
rect 55410 49758 55422 49810
rect 56466 49758 56478 49810
rect 56530 49758 56542 49810
rect 57486 49746 57538 49758
rect 57822 49810 57874 49822
rect 65326 49810 65378 49822
rect 61842 49758 61854 49810
rect 61906 49758 61918 49810
rect 62514 49758 62526 49810
rect 62578 49758 62590 49810
rect 57822 49746 57874 49758
rect 65326 49746 65378 49758
rect 66446 49810 66498 49822
rect 66446 49746 66498 49758
rect 68014 49810 68066 49822
rect 68014 49746 68066 49758
rect 69694 49810 69746 49822
rect 83022 49810 83074 49822
rect 86382 49810 86434 49822
rect 70354 49758 70366 49810
rect 70418 49758 70430 49810
rect 71250 49758 71262 49810
rect 71314 49758 71326 49810
rect 77522 49758 77534 49810
rect 77586 49758 77598 49810
rect 81778 49758 81790 49810
rect 81842 49758 81854 49810
rect 82226 49758 82238 49810
rect 82290 49758 82302 49810
rect 83570 49758 83582 49810
rect 83634 49758 83646 49810
rect 84354 49758 84366 49810
rect 84418 49758 84430 49810
rect 69694 49746 69746 49758
rect 83022 49746 83074 49758
rect 86382 49746 86434 49758
rect 86718 49810 86770 49822
rect 86718 49746 86770 49758
rect 87502 49810 87554 49822
rect 87502 49746 87554 49758
rect 87838 49810 87890 49822
rect 87838 49746 87890 49758
rect 88286 49810 88338 49822
rect 88286 49746 88338 49758
rect 89294 49810 89346 49822
rect 89294 49746 89346 49758
rect 89630 49810 89682 49822
rect 94558 49810 94610 49822
rect 94098 49758 94110 49810
rect 94162 49758 94174 49810
rect 89630 49746 89682 49758
rect 94558 49746 94610 49758
rect 97134 49810 97186 49822
rect 97134 49746 97186 49758
rect 97918 49810 97970 49822
rect 97918 49746 97970 49758
rect 58158 49698 58210 49710
rect 52546 49646 52558 49698
rect 52610 49646 52622 49698
rect 54674 49646 54686 49698
rect 54738 49646 54750 49698
rect 58158 49634 58210 49646
rect 58606 49698 58658 49710
rect 58606 49634 58658 49646
rect 61294 49698 61346 49710
rect 67454 49698 67506 49710
rect 81342 49698 81394 49710
rect 64642 49646 64654 49698
rect 64706 49646 64718 49698
rect 80434 49646 80446 49698
rect 80498 49646 80510 49698
rect 61294 49634 61346 49646
rect 67454 49634 67506 49646
rect 81342 49634 81394 49646
rect 85486 49698 85538 49710
rect 91186 49646 91198 49698
rect 91250 49646 91262 49698
rect 85486 49634 85538 49646
rect 66334 49586 66386 49598
rect 66334 49522 66386 49534
rect 88398 49586 88450 49598
rect 88398 49522 88450 49534
rect 90190 49586 90242 49598
rect 90190 49522 90242 49534
rect 1344 49418 98560 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 96638 49418
rect 96690 49366 96742 49418
rect 96794 49366 96846 49418
rect 96898 49366 98560 49418
rect 1344 49332 98560 49366
rect 54350 49250 54402 49262
rect 54350 49186 54402 49198
rect 61406 49138 61458 49150
rect 50530 49086 50542 49138
rect 50594 49086 50606 49138
rect 52658 49086 52670 49138
rect 52722 49086 52734 49138
rect 58706 49086 58718 49138
rect 58770 49086 58782 49138
rect 61406 49074 61458 49086
rect 76190 49138 76242 49150
rect 84366 49138 84418 49150
rect 79762 49086 79774 49138
rect 79826 49086 79838 49138
rect 81890 49086 81902 49138
rect 81954 49086 81966 49138
rect 76190 49074 76242 49086
rect 84366 49074 84418 49086
rect 86270 49138 86322 49150
rect 93214 49138 93266 49150
rect 88162 49086 88174 49138
rect 88226 49086 88238 49138
rect 94882 49086 94894 49138
rect 94946 49086 94958 49138
rect 97010 49086 97022 49138
rect 97074 49086 97086 49138
rect 86270 49074 86322 49086
rect 93214 49074 93266 49086
rect 68350 49026 68402 49038
rect 49858 48974 49870 49026
rect 49922 48974 49934 49026
rect 55794 48974 55806 49026
rect 55858 48974 55870 49026
rect 67106 48974 67118 49026
rect 67170 48974 67182 49026
rect 68350 48962 68402 48974
rect 68686 49026 68738 49038
rect 75742 49026 75794 49038
rect 69570 48974 69582 49026
rect 69634 48974 69646 49026
rect 68686 48962 68738 48974
rect 75742 48962 75794 48974
rect 77310 49026 77362 49038
rect 77310 48962 77362 48974
rect 78430 49026 78482 49038
rect 83918 49026 83970 49038
rect 79090 48974 79102 49026
rect 79154 48974 79166 49026
rect 78430 48962 78482 48974
rect 83918 48962 83970 48974
rect 85598 49026 85650 49038
rect 85598 48962 85650 48974
rect 85934 49026 85986 49038
rect 91970 48974 91982 49026
rect 92034 48974 92046 49026
rect 97682 48974 97694 49026
rect 97746 48974 97758 49026
rect 85934 48962 85986 48974
rect 53678 48914 53730 48926
rect 53678 48850 53730 48862
rect 54350 48914 54402 48926
rect 54350 48850 54402 48862
rect 54462 48914 54514 48926
rect 54462 48850 54514 48862
rect 55134 48914 55186 48926
rect 55134 48850 55186 48862
rect 55246 48914 55298 48926
rect 68462 48914 68514 48926
rect 77646 48914 77698 48926
rect 56578 48862 56590 48914
rect 56642 48862 56654 48914
rect 65202 48862 65214 48914
rect 65266 48862 65278 48914
rect 73154 48862 73166 48914
rect 73218 48862 73230 48914
rect 55246 48850 55298 48862
rect 68462 48850 68514 48862
rect 77646 48850 77698 48862
rect 83134 48914 83186 48926
rect 83134 48850 83186 48862
rect 83582 48914 83634 48926
rect 83582 48850 83634 48862
rect 83806 48914 83858 48926
rect 83806 48850 83858 48862
rect 85710 48914 85762 48926
rect 85710 48850 85762 48862
rect 93774 48914 93826 48926
rect 93774 48850 93826 48862
rect 94110 48914 94162 48926
rect 94110 48850 94162 48862
rect 53342 48802 53394 48814
rect 53342 48738 53394 48750
rect 53566 48802 53618 48814
rect 53566 48738 53618 48750
rect 54910 48802 54962 48814
rect 54910 48738 54962 48750
rect 60622 48802 60674 48814
rect 60622 48738 60674 48750
rect 67678 48802 67730 48814
rect 67678 48738 67730 48750
rect 75406 48802 75458 48814
rect 75406 48738 75458 48750
rect 78094 48802 78146 48814
rect 78094 48738 78146 48750
rect 78318 48802 78370 48814
rect 78318 48738 78370 48750
rect 82350 48802 82402 48814
rect 82350 48738 82402 48750
rect 82798 48802 82850 48814
rect 82798 48738 82850 48750
rect 83022 48802 83074 48814
rect 83022 48738 83074 48750
rect 1344 48634 98560 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 81278 48634
rect 81330 48582 81382 48634
rect 81434 48582 81486 48634
rect 81538 48582 98560 48634
rect 1344 48548 98560 48582
rect 53342 48466 53394 48478
rect 53342 48402 53394 48414
rect 53902 48466 53954 48478
rect 53902 48402 53954 48414
rect 57598 48466 57650 48478
rect 57598 48402 57650 48414
rect 58606 48466 58658 48478
rect 58606 48402 58658 48414
rect 61854 48466 61906 48478
rect 61854 48402 61906 48414
rect 62638 48466 62690 48478
rect 62638 48402 62690 48414
rect 63198 48466 63250 48478
rect 63198 48402 63250 48414
rect 64206 48466 64258 48478
rect 64206 48402 64258 48414
rect 67342 48466 67394 48478
rect 67342 48402 67394 48414
rect 68014 48466 68066 48478
rect 68014 48402 68066 48414
rect 72046 48466 72098 48478
rect 92654 48466 92706 48478
rect 78306 48414 78318 48466
rect 78370 48414 78382 48466
rect 72046 48402 72098 48414
rect 92654 48402 92706 48414
rect 97918 48466 97970 48478
rect 97918 48402 97970 48414
rect 53454 48354 53506 48366
rect 50530 48302 50542 48354
rect 50594 48302 50606 48354
rect 53454 48290 53506 48302
rect 54126 48354 54178 48366
rect 54126 48290 54178 48302
rect 54910 48354 54962 48366
rect 54910 48290 54962 48302
rect 55022 48354 55074 48366
rect 55022 48290 55074 48302
rect 56478 48354 56530 48366
rect 56478 48290 56530 48302
rect 57374 48354 57426 48366
rect 57374 48290 57426 48302
rect 58270 48354 58322 48366
rect 58270 48290 58322 48302
rect 58382 48354 58434 48366
rect 58382 48290 58434 48302
rect 59166 48354 59218 48366
rect 59166 48290 59218 48302
rect 60734 48354 60786 48366
rect 60734 48290 60786 48302
rect 62526 48354 62578 48366
rect 62526 48290 62578 48302
rect 62862 48354 62914 48366
rect 62862 48290 62914 48302
rect 63422 48354 63474 48366
rect 63422 48290 63474 48302
rect 63534 48354 63586 48366
rect 63534 48290 63586 48302
rect 65550 48354 65602 48366
rect 65550 48290 65602 48302
rect 66334 48354 66386 48366
rect 72270 48354 72322 48366
rect 69458 48302 69470 48354
rect 69522 48302 69534 48354
rect 66334 48290 66386 48302
rect 72270 48290 72322 48302
rect 72382 48354 72434 48366
rect 72382 48290 72434 48302
rect 78766 48354 78818 48366
rect 92878 48354 92930 48366
rect 82338 48302 82350 48354
rect 82402 48302 82414 48354
rect 87154 48302 87166 48354
rect 87218 48302 87230 48354
rect 90066 48302 90078 48354
rect 90130 48302 90142 48354
rect 78766 48290 78818 48302
rect 92878 48290 92930 48302
rect 92990 48354 93042 48366
rect 92990 48290 93042 48302
rect 97358 48354 97410 48366
rect 97358 48290 97410 48302
rect 97470 48354 97522 48366
rect 97470 48290 97522 48302
rect 53118 48242 53170 48254
rect 49858 48190 49870 48242
rect 49922 48190 49934 48242
rect 53118 48178 53170 48190
rect 54238 48242 54290 48254
rect 54238 48178 54290 48190
rect 56254 48242 56306 48254
rect 56254 48178 56306 48190
rect 56590 48242 56642 48254
rect 56590 48178 56642 48190
rect 57710 48242 57762 48254
rect 57710 48178 57762 48190
rect 58942 48242 58994 48254
rect 58942 48178 58994 48190
rect 59278 48242 59330 48254
rect 59278 48178 59330 48190
rect 60622 48242 60674 48254
rect 60622 48178 60674 48190
rect 60958 48242 61010 48254
rect 60958 48178 61010 48190
rect 61966 48242 62018 48254
rect 61966 48178 62018 48190
rect 64318 48242 64370 48254
rect 64318 48178 64370 48190
rect 65326 48242 65378 48254
rect 65326 48178 65378 48190
rect 65662 48242 65714 48254
rect 65662 48178 65714 48190
rect 66110 48242 66162 48254
rect 66110 48178 66162 48190
rect 66446 48242 66498 48254
rect 66446 48178 66498 48190
rect 67902 48242 67954 48254
rect 67902 48178 67954 48190
rect 68238 48242 68290 48254
rect 68674 48190 68686 48242
rect 68738 48190 68750 48242
rect 76738 48190 76750 48242
rect 76802 48190 76814 48242
rect 77634 48190 77646 48242
rect 77698 48190 77710 48242
rect 78082 48190 78094 48242
rect 78146 48190 78158 48242
rect 79538 48190 79550 48242
rect 79602 48190 79614 48242
rect 80434 48190 80446 48242
rect 80498 48190 80510 48242
rect 81666 48190 81678 48242
rect 81730 48190 81742 48242
rect 87938 48190 87950 48242
rect 88002 48190 88014 48242
rect 89282 48190 89294 48242
rect 89346 48190 89358 48242
rect 93650 48190 93662 48242
rect 93714 48190 93726 48242
rect 68238 48178 68290 48190
rect 55470 48130 55522 48142
rect 52658 48078 52670 48130
rect 52722 48078 52734 48130
rect 55470 48066 55522 48078
rect 59726 48130 59778 48142
rect 59726 48066 59778 48078
rect 66894 48130 66946 48142
rect 73278 48130 73330 48142
rect 77310 48130 77362 48142
rect 88622 48130 88674 48142
rect 71586 48078 71598 48130
rect 71650 48078 71662 48130
rect 73826 48078 73838 48130
rect 73890 48078 73902 48130
rect 75954 48078 75966 48130
rect 76018 48078 76030 48130
rect 84466 48078 84478 48130
rect 84530 48078 84542 48130
rect 85026 48078 85038 48130
rect 85090 48078 85102 48130
rect 92194 48078 92206 48130
rect 92258 48078 92270 48130
rect 94322 48078 94334 48130
rect 94386 48078 94398 48130
rect 96450 48078 96462 48130
rect 96514 48078 96526 48130
rect 66894 48066 66946 48078
rect 73278 48066 73330 48078
rect 77310 48066 77362 48078
rect 88622 48066 88674 48078
rect 54910 48018 54962 48030
rect 54910 47954 54962 47966
rect 61854 48018 61906 48030
rect 61854 47954 61906 47966
rect 64206 48018 64258 48030
rect 64206 47954 64258 47966
rect 97358 48018 97410 48030
rect 97358 47954 97410 47966
rect 1344 47850 98560 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 96638 47850
rect 96690 47798 96742 47850
rect 96794 47798 96846 47850
rect 96898 47798 98560 47850
rect 1344 47764 98560 47798
rect 59950 47570 60002 47582
rect 50082 47518 50094 47570
rect 50146 47518 50158 47570
rect 52210 47518 52222 47570
rect 52274 47518 52286 47570
rect 55794 47518 55806 47570
rect 55858 47518 55870 47570
rect 59950 47506 60002 47518
rect 60622 47570 60674 47582
rect 60622 47506 60674 47518
rect 62078 47570 62130 47582
rect 67006 47570 67058 47582
rect 62850 47518 62862 47570
rect 62914 47518 62926 47570
rect 62078 47506 62130 47518
rect 67006 47506 67058 47518
rect 67790 47570 67842 47582
rect 67790 47506 67842 47518
rect 70814 47570 70866 47582
rect 76414 47570 76466 47582
rect 75842 47518 75854 47570
rect 75906 47518 75918 47570
rect 70814 47506 70866 47518
rect 76414 47506 76466 47518
rect 78654 47570 78706 47582
rect 78654 47506 78706 47518
rect 81006 47570 81058 47582
rect 81006 47506 81058 47518
rect 82238 47570 82290 47582
rect 82238 47506 82290 47518
rect 83470 47570 83522 47582
rect 83470 47506 83522 47518
rect 84142 47570 84194 47582
rect 84142 47506 84194 47518
rect 84478 47570 84530 47582
rect 94782 47570 94834 47582
rect 89954 47518 89966 47570
rect 90018 47518 90030 47570
rect 92082 47518 92094 47570
rect 92146 47518 92158 47570
rect 84478 47506 84530 47518
rect 94782 47506 94834 47518
rect 97246 47570 97298 47582
rect 97246 47506 97298 47518
rect 61742 47458 61794 47470
rect 66558 47458 66610 47470
rect 49410 47406 49422 47458
rect 49474 47406 49486 47458
rect 54898 47406 54910 47458
rect 54962 47406 54974 47458
rect 65762 47406 65774 47458
rect 65826 47406 65838 47458
rect 61742 47394 61794 47406
rect 66558 47394 66610 47406
rect 69582 47458 69634 47470
rect 69582 47394 69634 47406
rect 72158 47458 72210 47470
rect 73042 47418 73054 47470
rect 73106 47418 73118 47470
rect 77198 47458 77250 47470
rect 86942 47458 86994 47470
rect 96126 47458 96178 47470
rect 72158 47394 72210 47406
rect 85586 47406 85598 47458
rect 85650 47406 85662 47458
rect 86482 47406 86494 47458
rect 86546 47406 86558 47458
rect 87714 47406 87726 47458
rect 87778 47406 87790 47458
rect 88162 47406 88174 47458
rect 88226 47406 88238 47458
rect 89282 47406 89294 47458
rect 89346 47406 89358 47458
rect 77198 47394 77250 47406
rect 86942 47394 86994 47406
rect 96126 47394 96178 47406
rect 96462 47458 96514 47470
rect 96462 47394 96514 47406
rect 61406 47346 61458 47358
rect 61406 47282 61458 47294
rect 61518 47346 61570 47358
rect 68462 47346 68514 47358
rect 64978 47294 64990 47346
rect 65042 47294 65054 47346
rect 61518 47282 61570 47294
rect 68462 47282 68514 47294
rect 68574 47346 68626 47358
rect 68574 47282 68626 47294
rect 69470 47346 69522 47358
rect 69470 47282 69522 47294
rect 70030 47346 70082 47358
rect 70030 47282 70082 47294
rect 70366 47346 70418 47358
rect 70366 47282 70418 47294
rect 72270 47346 72322 47358
rect 78206 47346 78258 47358
rect 73714 47294 73726 47346
rect 73778 47294 73790 47346
rect 72270 47282 72322 47294
rect 78206 47282 78258 47294
rect 88622 47346 88674 47358
rect 88622 47282 88674 47294
rect 93214 47346 93266 47358
rect 93214 47282 93266 47294
rect 93550 47346 93602 47358
rect 93550 47282 93602 47294
rect 94334 47346 94386 47358
rect 94334 47282 94386 47294
rect 95230 47346 95282 47358
rect 95230 47282 95282 47294
rect 96238 47346 96290 47358
rect 96238 47282 96290 47294
rect 52670 47234 52722 47246
rect 52670 47170 52722 47182
rect 59502 47234 59554 47246
rect 59502 47170 59554 47182
rect 66222 47234 66274 47246
rect 66222 47170 66274 47182
rect 66446 47234 66498 47246
rect 66446 47170 66498 47182
rect 68238 47234 68290 47246
rect 68238 47170 68290 47182
rect 69246 47234 69298 47246
rect 69246 47170 69298 47182
rect 70254 47234 70306 47246
rect 70254 47170 70306 47182
rect 71262 47234 71314 47246
rect 71262 47170 71314 47182
rect 72494 47234 72546 47246
rect 72494 47170 72546 47182
rect 77646 47234 77698 47246
rect 93998 47234 94050 47246
rect 87602 47182 87614 47234
rect 87666 47182 87678 47234
rect 77646 47170 77698 47182
rect 93998 47170 94050 47182
rect 94222 47234 94274 47246
rect 94222 47170 94274 47182
rect 96798 47234 96850 47246
rect 96798 47170 96850 47182
rect 1344 47066 98560 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 81278 47066
rect 81330 47014 81382 47066
rect 81434 47014 81486 47066
rect 81538 47014 98560 47066
rect 1344 46980 98560 47014
rect 53342 46898 53394 46910
rect 53342 46834 53394 46846
rect 53566 46898 53618 46910
rect 53566 46834 53618 46846
rect 54238 46898 54290 46910
rect 54238 46834 54290 46846
rect 55246 46898 55298 46910
rect 55246 46834 55298 46846
rect 55694 46898 55746 46910
rect 55694 46834 55746 46846
rect 56030 46898 56082 46910
rect 56030 46834 56082 46846
rect 57486 46898 57538 46910
rect 57486 46834 57538 46846
rect 66222 46898 66274 46910
rect 66222 46834 66274 46846
rect 70590 46898 70642 46910
rect 70590 46834 70642 46846
rect 71934 46898 71986 46910
rect 71934 46834 71986 46846
rect 72718 46898 72770 46910
rect 72718 46834 72770 46846
rect 73278 46898 73330 46910
rect 73278 46834 73330 46846
rect 73950 46898 74002 46910
rect 73950 46834 74002 46846
rect 75630 46898 75682 46910
rect 75630 46834 75682 46846
rect 75854 46898 75906 46910
rect 75854 46834 75906 46846
rect 76414 46898 76466 46910
rect 76414 46834 76466 46846
rect 77534 46898 77586 46910
rect 77534 46834 77586 46846
rect 77982 46898 78034 46910
rect 77982 46834 78034 46846
rect 82462 46898 82514 46910
rect 82462 46834 82514 46846
rect 85150 46898 85202 46910
rect 85150 46834 85202 46846
rect 93214 46898 93266 46910
rect 93214 46834 93266 46846
rect 93438 46898 93490 46910
rect 93438 46834 93490 46846
rect 93774 46898 93826 46910
rect 93774 46834 93826 46846
rect 95118 46898 95170 46910
rect 95118 46834 95170 46846
rect 95678 46898 95730 46910
rect 95678 46834 95730 46846
rect 96014 46898 96066 46910
rect 96014 46834 96066 46846
rect 96574 46898 96626 46910
rect 96574 46834 96626 46846
rect 53678 46786 53730 46798
rect 65550 46786 65602 46798
rect 62178 46734 62190 46786
rect 62242 46734 62254 46786
rect 53678 46722 53730 46734
rect 65550 46722 65602 46734
rect 65662 46786 65714 46798
rect 65662 46722 65714 46734
rect 73838 46786 73890 46798
rect 73838 46722 73890 46734
rect 75070 46786 75122 46798
rect 75070 46722 75122 46734
rect 75518 46786 75570 46798
rect 75518 46722 75570 46734
rect 76302 46786 76354 46798
rect 93102 46786 93154 46798
rect 87714 46734 87726 46786
rect 87778 46734 87790 46786
rect 76302 46722 76354 46734
rect 93102 46722 93154 46734
rect 61506 46622 61518 46674
rect 61570 46622 61582 46674
rect 66882 46622 66894 46674
rect 66946 46622 66958 46674
rect 82226 46622 82238 46674
rect 82290 46622 82302 46674
rect 88386 46622 88398 46674
rect 88450 46622 88462 46674
rect 89618 46622 89630 46674
rect 89682 46622 89694 46674
rect 52446 46562 52498 46574
rect 52446 46498 52498 46510
rect 52894 46562 52946 46574
rect 52894 46498 52946 46510
rect 54798 46562 54850 46574
rect 54798 46498 54850 46510
rect 60958 46562 61010 46574
rect 70142 46562 70194 46574
rect 64306 46510 64318 46562
rect 64370 46510 64382 46562
rect 67554 46510 67566 46562
rect 67618 46510 67630 46562
rect 69682 46510 69694 46562
rect 69746 46510 69758 46562
rect 60958 46498 61010 46510
rect 70142 46498 70194 46510
rect 76974 46562 77026 46574
rect 76974 46498 77026 46510
rect 81678 46562 81730 46574
rect 94334 46562 94386 46574
rect 85586 46510 85598 46562
rect 85650 46510 85662 46562
rect 90402 46510 90414 46562
rect 90466 46510 90478 46562
rect 92530 46510 92542 46562
rect 92594 46510 92606 46562
rect 81678 46498 81730 46510
rect 94334 46498 94386 46510
rect 94782 46562 94834 46574
rect 94782 46498 94834 46510
rect 65550 46450 65602 46462
rect 54450 46398 54462 46450
rect 54514 46447 54526 46450
rect 54786 46447 54798 46450
rect 54514 46401 54798 46447
rect 54514 46398 54526 46401
rect 54786 46398 54798 46401
rect 54850 46398 54862 46450
rect 55458 46398 55470 46450
rect 55522 46447 55534 46450
rect 56018 46447 56030 46450
rect 55522 46401 56030 46447
rect 55522 46398 55534 46401
rect 56018 46398 56030 46401
rect 56082 46398 56094 46450
rect 65550 46386 65602 46398
rect 73950 46450 74002 46462
rect 73950 46386 74002 46398
rect 76414 46450 76466 46462
rect 94770 46398 94782 46450
rect 94834 46447 94846 46450
rect 95666 46447 95678 46450
rect 94834 46401 95678 46447
rect 94834 46398 94846 46401
rect 95666 46398 95678 46401
rect 95730 46398 95742 46450
rect 76414 46386 76466 46398
rect 1344 46282 98560 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 98560 46282
rect 1344 46196 98560 46230
rect 64990 46114 65042 46126
rect 94322 46062 94334 46114
rect 94386 46111 94398 46114
rect 95330 46111 95342 46114
rect 94386 46065 95342 46111
rect 94386 46062 94398 46065
rect 95330 46062 95342 46065
rect 95394 46062 95406 46114
rect 64990 46050 65042 46062
rect 75294 46002 75346 46014
rect 56130 45950 56142 46002
rect 56194 45950 56206 46002
rect 58258 45950 58270 46002
rect 58322 45950 58334 46002
rect 62178 45950 62190 46002
rect 62242 45950 62254 46002
rect 64306 45950 64318 46002
rect 64370 45950 64382 46002
rect 75294 45938 75346 45950
rect 76078 46002 76130 46014
rect 76078 45938 76130 45950
rect 83918 46002 83970 46014
rect 83918 45938 83970 45950
rect 89070 46002 89122 46014
rect 89070 45938 89122 45950
rect 91310 46002 91362 46014
rect 91310 45938 91362 45950
rect 92430 46002 92482 46014
rect 92430 45938 92482 45950
rect 94110 46002 94162 46014
rect 94110 45938 94162 45950
rect 94670 46002 94722 46014
rect 94670 45938 94722 45950
rect 95118 46002 95170 46014
rect 95118 45938 95170 45950
rect 65102 45890 65154 45902
rect 55458 45838 55470 45890
rect 55522 45838 55534 45890
rect 61506 45838 61518 45890
rect 61570 45838 61582 45890
rect 65102 45826 65154 45838
rect 68126 45890 68178 45902
rect 68126 45826 68178 45838
rect 68462 45890 68514 45902
rect 82238 45890 82290 45902
rect 81330 45838 81342 45890
rect 81394 45838 81406 45890
rect 68462 45826 68514 45838
rect 82238 45826 82290 45838
rect 82574 45890 82626 45902
rect 82574 45826 82626 45838
rect 85710 45890 85762 45902
rect 85710 45826 85762 45838
rect 89742 45890 89794 45902
rect 89742 45826 89794 45838
rect 90078 45890 90130 45902
rect 90078 45826 90130 45838
rect 90526 45890 90578 45902
rect 90526 45826 90578 45838
rect 90862 45890 90914 45902
rect 90862 45826 90914 45838
rect 51214 45778 51266 45790
rect 51214 45714 51266 45726
rect 64990 45778 65042 45790
rect 64990 45714 65042 45726
rect 68350 45778 68402 45790
rect 68350 45714 68402 45726
rect 79102 45778 79154 45790
rect 79102 45714 79154 45726
rect 80670 45778 80722 45790
rect 84478 45778 84530 45790
rect 89854 45778 89906 45790
rect 82786 45726 82798 45778
rect 82850 45726 82862 45778
rect 83122 45726 83134 45778
rect 83186 45726 83198 45778
rect 85922 45726 85934 45778
rect 85986 45726 85998 45778
rect 86258 45726 86270 45778
rect 86322 45726 86334 45778
rect 80670 45714 80722 45726
rect 84478 45714 84530 45726
rect 89854 45714 89906 45726
rect 90750 45778 90802 45790
rect 90750 45714 90802 45726
rect 50878 45666 50930 45678
rect 50878 45602 50930 45614
rect 58718 45666 58770 45678
rect 58718 45602 58770 45614
rect 70142 45666 70194 45678
rect 70142 45602 70194 45614
rect 77310 45666 77362 45678
rect 77310 45602 77362 45614
rect 78766 45666 78818 45678
rect 78766 45602 78818 45614
rect 81566 45666 81618 45678
rect 81566 45602 81618 45614
rect 85374 45666 85426 45678
rect 85374 45602 85426 45614
rect 91982 45666 92034 45678
rect 91982 45602 92034 45614
rect 93102 45666 93154 45678
rect 93102 45602 93154 45614
rect 93550 45666 93602 45678
rect 93550 45602 93602 45614
rect 95566 45666 95618 45678
rect 95566 45602 95618 45614
rect 95902 45666 95954 45678
rect 95902 45602 95954 45614
rect 1344 45498 98560 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 98560 45498
rect 1344 45412 98560 45446
rect 70926 45330 70978 45342
rect 70926 45266 70978 45278
rect 71374 45330 71426 45342
rect 75070 45330 75122 45342
rect 74722 45278 74734 45330
rect 74786 45278 74798 45330
rect 71374 45266 71426 45278
rect 75070 45266 75122 45278
rect 56254 45218 56306 45230
rect 75630 45218 75682 45230
rect 50754 45166 50766 45218
rect 50818 45166 50830 45218
rect 63522 45166 63534 45218
rect 63586 45166 63598 45218
rect 67666 45166 67678 45218
rect 67730 45166 67742 45218
rect 56254 45154 56306 45166
rect 75630 45154 75682 45166
rect 77086 45218 77138 45230
rect 96126 45218 96178 45230
rect 78418 45166 78430 45218
rect 78482 45166 78494 45218
rect 82114 45166 82126 45218
rect 82178 45166 82190 45218
rect 91970 45166 91982 45218
rect 92034 45166 92046 45218
rect 77086 45154 77138 45166
rect 96126 45154 96178 45166
rect 56590 45106 56642 45118
rect 75966 45106 76018 45118
rect 50082 45054 50094 45106
rect 50146 45054 50158 45106
rect 64194 45054 64206 45106
rect 64258 45054 64270 45106
rect 66994 45054 67006 45106
rect 67058 45054 67070 45106
rect 56590 45042 56642 45054
rect 75966 45042 76018 45054
rect 76750 45106 76802 45118
rect 95790 45106 95842 45118
rect 77746 45054 77758 45106
rect 77810 45054 77822 45106
rect 81330 45054 81342 45106
rect 81394 45054 81406 45106
rect 84914 45054 84926 45106
rect 84978 45054 84990 45106
rect 91410 45054 91422 45106
rect 91474 45054 91486 45106
rect 76750 45042 76802 45054
rect 95790 45042 95842 45054
rect 53454 44994 53506 45006
rect 70366 44994 70418 45006
rect 88174 44994 88226 45006
rect 52882 44942 52894 44994
rect 52946 44942 52958 44994
rect 61394 44942 61406 44994
rect 61458 44942 61470 44994
rect 69794 44942 69806 44994
rect 69858 44942 69870 44994
rect 80546 44942 80558 44994
rect 80610 44942 80622 44994
rect 84242 44942 84254 44994
rect 84306 44942 84318 44994
rect 85586 44942 85598 44994
rect 85650 44942 85662 44994
rect 87714 44942 87726 44994
rect 87778 44942 87790 44994
rect 53454 44930 53506 44942
rect 70366 44930 70418 44942
rect 88174 44930 88226 44942
rect 1344 44714 98560 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 98560 44714
rect 1344 44628 98560 44662
rect 77422 44546 77474 44558
rect 93314 44494 93326 44546
rect 93378 44543 93390 44546
rect 93986 44543 93998 44546
rect 93378 44497 93998 44543
rect 93378 44494 93390 44497
rect 93986 44494 93998 44497
rect 94050 44494 94062 44546
rect 77422 44482 77474 44494
rect 58606 44434 58658 44446
rect 51874 44382 51886 44434
rect 51938 44382 51950 44434
rect 56018 44382 56030 44434
rect 56082 44382 56094 44434
rect 58146 44382 58158 44434
rect 58210 44382 58222 44434
rect 58606 44370 58658 44382
rect 59278 44434 59330 44446
rect 59278 44370 59330 44382
rect 61854 44434 61906 44446
rect 77758 44434 77810 44446
rect 93102 44434 93154 44446
rect 72370 44382 72382 44434
rect 72434 44382 72446 44434
rect 74386 44382 74398 44434
rect 74450 44382 74462 44434
rect 76514 44382 76526 44434
rect 76578 44382 76590 44434
rect 80658 44382 80670 44434
rect 80722 44382 80734 44434
rect 61854 44370 61906 44382
rect 77758 44370 77810 44382
rect 93102 44370 93154 44382
rect 93998 44434 94050 44446
rect 94882 44382 94894 44434
rect 94946 44382 94958 44434
rect 97010 44382 97022 44434
rect 97074 44382 97086 44434
rect 93998 44370 94050 44382
rect 91982 44322 92034 44334
rect 49074 44270 49086 44322
rect 49138 44270 49150 44322
rect 55346 44270 55358 44322
rect 55410 44270 55422 44322
rect 62514 44270 62526 44322
rect 62578 44270 62590 44322
rect 67218 44270 67230 44322
rect 67282 44270 67294 44322
rect 69458 44270 69470 44322
rect 69522 44270 69534 44322
rect 73714 44270 73726 44322
rect 73778 44270 73790 44322
rect 83906 44270 83918 44322
rect 83970 44270 83982 44322
rect 85362 44270 85374 44322
rect 85426 44270 85438 44322
rect 91298 44270 91310 44322
rect 91362 44270 91374 44322
rect 91982 44258 92034 44270
rect 93550 44322 93602 44334
rect 97682 44270 97694 44322
rect 97746 44270 97758 44322
rect 93550 44258 93602 44270
rect 85598 44210 85650 44222
rect 49746 44158 49758 44210
rect 49810 44158 49822 44210
rect 66322 44158 66334 44210
rect 66386 44158 66398 44210
rect 70242 44158 70254 44210
rect 70306 44158 70318 44210
rect 77970 44158 77982 44210
rect 78034 44158 78046 44210
rect 78530 44158 78542 44210
rect 78594 44158 78606 44210
rect 91186 44158 91198 44210
rect 91250 44158 91262 44210
rect 85598 44146 85650 44158
rect 52334 44098 52386 44110
rect 52334 44034 52386 44046
rect 62750 44098 62802 44110
rect 62750 44034 62802 44046
rect 72830 44098 72882 44110
rect 72830 44034 72882 44046
rect 90638 44098 90690 44110
rect 90638 44034 90690 44046
rect 92318 44098 92370 44110
rect 92318 44034 92370 44046
rect 1344 43930 98560 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 98560 43930
rect 1344 43844 98560 43878
rect 48750 43762 48802 43774
rect 48750 43698 48802 43710
rect 63422 43762 63474 43774
rect 63422 43698 63474 43710
rect 70254 43762 70306 43774
rect 70254 43698 70306 43710
rect 76302 43762 76354 43774
rect 76302 43698 76354 43710
rect 51662 43650 51714 43662
rect 54350 43650 54402 43662
rect 50754 43598 50766 43650
rect 50818 43598 50830 43650
rect 52210 43598 52222 43650
rect 52274 43598 52286 43650
rect 52770 43598 52782 43650
rect 52834 43598 52846 43650
rect 51662 43586 51714 43598
rect 54350 43586 54402 43598
rect 55022 43650 55074 43662
rect 55022 43586 55074 43598
rect 56702 43650 56754 43662
rect 56702 43586 56754 43598
rect 57598 43650 57650 43662
rect 59838 43650 59890 43662
rect 72718 43650 72770 43662
rect 97134 43650 97186 43662
rect 58482 43598 58494 43650
rect 58546 43598 58558 43650
rect 64418 43598 64430 43650
rect 64482 43598 64494 43650
rect 71474 43598 71486 43650
rect 71538 43598 71550 43650
rect 72034 43598 72046 43650
rect 72098 43598 72110 43650
rect 75282 43598 75294 43650
rect 75346 43598 75358 43650
rect 77858 43598 77870 43650
rect 77922 43598 77934 43650
rect 95554 43598 95566 43650
rect 95618 43598 95630 43650
rect 57598 43586 57650 43598
rect 59838 43586 59890 43598
rect 72718 43586 72770 43598
rect 97134 43586 97186 43598
rect 49758 43538 49810 43550
rect 53790 43538 53842 43550
rect 48514 43486 48526 43538
rect 48578 43486 48590 43538
rect 50866 43486 50878 43538
rect 50930 43486 50942 43538
rect 49758 43474 49810 43486
rect 53790 43474 53842 43486
rect 55358 43538 55410 43550
rect 60174 43538 60226 43550
rect 65774 43538 65826 43550
rect 70926 43538 70978 43550
rect 58706 43486 58718 43538
rect 58770 43486 58782 43538
rect 64530 43486 64542 43538
rect 64594 43486 64606 43538
rect 70018 43486 70030 43538
rect 70082 43486 70094 43538
rect 55358 43474 55410 43486
rect 60174 43474 60226 43486
rect 65774 43474 65826 43486
rect 70926 43474 70978 43486
rect 71262 43538 71314 43550
rect 71262 43474 71314 43486
rect 74622 43538 74674 43550
rect 75966 43538 76018 43550
rect 75170 43486 75182 43538
rect 75234 43486 75246 43538
rect 77186 43486 77198 43538
rect 77250 43486 77262 43538
rect 92642 43486 92654 43538
rect 92706 43486 92718 43538
rect 74622 43474 74674 43486
rect 75966 43474 76018 43486
rect 50094 43426 50146 43438
rect 50094 43362 50146 43374
rect 51998 43426 52050 43438
rect 51998 43362 52050 43374
rect 53342 43426 53394 43438
rect 53342 43362 53394 43374
rect 59278 43426 59330 43438
rect 59278 43362 59330 43374
rect 65326 43426 65378 43438
rect 65326 43362 65378 43374
rect 69358 43426 69410 43438
rect 84702 43426 84754 43438
rect 79986 43374 79998 43426
rect 80050 43374 80062 43426
rect 69358 43362 69410 43374
rect 84702 43362 84754 43374
rect 89742 43426 89794 43438
rect 89742 43362 89794 43374
rect 90078 43426 90130 43438
rect 90078 43362 90130 43374
rect 57934 43314 57986 43326
rect 57934 43250 57986 43262
rect 63758 43314 63810 43326
rect 63758 43250 63810 43262
rect 1344 43146 98560 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 98560 43146
rect 1344 43060 98560 43094
rect 77422 42978 77474 42990
rect 77422 42914 77474 42926
rect 77758 42978 77810 42990
rect 77758 42914 77810 42926
rect 53454 42866 53506 42878
rect 62526 42866 62578 42878
rect 68574 42866 68626 42878
rect 79214 42866 79266 42878
rect 52658 42814 52670 42866
rect 52722 42814 52734 42866
rect 54786 42814 54798 42866
rect 54850 42814 54862 42866
rect 56914 42814 56926 42866
rect 56978 42814 56990 42866
rect 60386 42814 60398 42866
rect 60450 42814 60462 42866
rect 63858 42814 63870 42866
rect 63922 42814 63934 42866
rect 65986 42814 65998 42866
rect 66050 42814 66062 42866
rect 72258 42814 72270 42866
rect 72322 42814 72334 42866
rect 53454 42802 53506 42814
rect 62526 42802 62578 42814
rect 68574 42802 68626 42814
rect 79214 42802 79266 42814
rect 87502 42866 87554 42878
rect 87502 42802 87554 42814
rect 94334 42866 94386 42878
rect 94882 42814 94894 42866
rect 94946 42814 94958 42866
rect 94334 42802 94386 42814
rect 75742 42754 75794 42766
rect 86158 42754 86210 42766
rect 49746 42702 49758 42754
rect 49810 42702 49822 42754
rect 54114 42702 54126 42754
rect 54178 42702 54190 42754
rect 57586 42702 57598 42754
rect 57650 42702 57662 42754
rect 63074 42702 63086 42754
rect 63138 42702 63150 42754
rect 69346 42702 69358 42754
rect 69410 42702 69422 42754
rect 81778 42702 81790 42754
rect 81842 42702 81854 42754
rect 75742 42690 75794 42702
rect 86158 42690 86210 42702
rect 89742 42754 89794 42766
rect 89742 42690 89794 42702
rect 93214 42754 93266 42766
rect 97682 42702 97694 42754
rect 97746 42702 97758 42754
rect 93214 42690 93266 42702
rect 85262 42642 85314 42654
rect 50530 42590 50542 42642
rect 50594 42590 50606 42642
rect 58258 42590 58270 42642
rect 58322 42590 58334 42642
rect 77970 42590 77982 42642
rect 78034 42590 78046 42642
rect 78530 42590 78542 42642
rect 78594 42590 78606 42642
rect 86370 42590 86382 42642
rect 86434 42590 86446 42642
rect 86930 42590 86942 42642
rect 86994 42590 87006 42642
rect 89954 42590 89966 42642
rect 90018 42590 90030 42642
rect 90514 42590 90526 42642
rect 90578 42590 90590 42642
rect 97010 42590 97022 42642
rect 97074 42590 97086 42642
rect 85262 42578 85314 42590
rect 61294 42530 61346 42542
rect 61294 42466 61346 42478
rect 62078 42530 62130 42542
rect 62078 42466 62130 42478
rect 66446 42530 66498 42542
rect 66446 42466 66498 42478
rect 75182 42530 75234 42542
rect 75182 42466 75234 42478
rect 76190 42530 76242 42542
rect 76190 42466 76242 42478
rect 82014 42530 82066 42542
rect 82014 42466 82066 42478
rect 85822 42530 85874 42542
rect 85822 42466 85874 42478
rect 88286 42530 88338 42542
rect 88286 42466 88338 42478
rect 88734 42530 88786 42542
rect 88734 42466 88786 42478
rect 89406 42530 89458 42542
rect 89406 42466 89458 42478
rect 92430 42530 92482 42542
rect 92430 42466 92482 42478
rect 93550 42530 93602 42542
rect 93550 42466 93602 42478
rect 1344 42362 98560 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 98560 42362
rect 1344 42276 98560 42310
rect 54798 42194 54850 42206
rect 54798 42130 54850 42142
rect 71710 42194 71762 42206
rect 71710 42130 71762 42142
rect 77758 42194 77810 42206
rect 77758 42130 77810 42142
rect 97246 42194 97298 42206
rect 97246 42130 97298 42142
rect 65438 42082 65490 42094
rect 54114 42030 54126 42082
rect 54178 42030 54190 42082
rect 56578 42030 56590 42082
rect 56642 42030 56654 42082
rect 60722 42030 60734 42082
rect 60786 42030 60798 42082
rect 64306 42030 64318 42082
rect 64370 42030 64382 42082
rect 65438 42018 65490 42030
rect 65774 42082 65826 42094
rect 70802 42030 70814 42082
rect 70866 42030 70878 42082
rect 82114 42030 82126 42082
rect 82178 42030 82190 42082
rect 95330 42030 95342 42082
rect 95394 42030 95406 42082
rect 65774 42018 65826 42030
rect 55470 41970 55522 41982
rect 73278 41970 73330 41982
rect 88174 41970 88226 41982
rect 96350 41970 96402 41982
rect 98030 41970 98082 41982
rect 49634 41918 49646 41970
rect 49698 41918 49710 41970
rect 54226 41918 54238 41970
rect 54290 41918 54302 41970
rect 56466 41918 56478 41970
rect 56530 41918 56542 41970
rect 62066 41918 62078 41970
rect 62130 41918 62142 41970
rect 64418 41918 64430 41970
rect 64482 41918 64494 41970
rect 66322 41918 66334 41970
rect 66386 41918 66398 41970
rect 70914 41918 70926 41970
rect 70978 41918 70990 41970
rect 73938 41918 73950 41970
rect 74002 41918 74014 41970
rect 81330 41918 81342 41970
rect 81394 41918 81406 41970
rect 84914 41918 84926 41970
rect 84978 41918 84990 41970
rect 89282 41918 89294 41970
rect 89346 41918 89358 41970
rect 95218 41918 95230 41970
rect 95282 41918 95294 41970
rect 97458 41918 97470 41970
rect 97522 41918 97534 41970
rect 55470 41906 55522 41918
rect 73278 41906 73330 41918
rect 88174 41906 88226 41918
rect 96350 41906 96402 41918
rect 98030 41906 98082 41918
rect 53454 41858 53506 41870
rect 50306 41806 50318 41858
rect 50370 41806 50382 41858
rect 52434 41806 52446 41858
rect 52498 41806 52510 41858
rect 53454 41794 53506 41806
rect 63422 41858 63474 41870
rect 77310 41858 77362 41870
rect 67106 41806 67118 41858
rect 67170 41806 67182 41858
rect 69234 41806 69246 41858
rect 69298 41806 69310 41858
rect 72146 41806 72158 41858
rect 72210 41806 72222 41858
rect 74722 41806 74734 41858
rect 74786 41806 74798 41858
rect 76850 41806 76862 41858
rect 76914 41806 76926 41858
rect 63422 41794 63474 41806
rect 77310 41794 77362 41806
rect 78206 41858 78258 41870
rect 84242 41806 84254 41858
rect 84306 41806 84318 41858
rect 85586 41806 85598 41858
rect 85650 41806 85662 41858
rect 87714 41806 87726 41858
rect 87778 41806 87790 41858
rect 94322 41806 94334 41858
rect 94386 41806 94398 41858
rect 78206 41794 78258 41806
rect 53118 41746 53170 41758
rect 53118 41682 53170 41694
rect 55806 41746 55858 41758
rect 55806 41682 55858 41694
rect 63758 41746 63810 41758
rect 63758 41682 63810 41694
rect 69918 41746 69970 41758
rect 69918 41682 69970 41694
rect 70254 41746 70306 41758
rect 70254 41682 70306 41694
rect 96014 41746 96066 41758
rect 96014 41682 96066 41694
rect 1344 41578 98560 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 98560 41578
rect 1344 41492 98560 41526
rect 51774 41410 51826 41422
rect 58942 41410 58994 41422
rect 53218 41358 53230 41410
rect 53282 41407 53294 41410
rect 53778 41407 53790 41410
rect 53282 41361 53790 41407
rect 53282 41358 53294 41361
rect 53778 41358 53790 41361
rect 53842 41358 53854 41410
rect 51774 41346 51826 41358
rect 58942 41346 58994 41358
rect 82126 41410 82178 41422
rect 82126 41346 82178 41358
rect 90302 41410 90354 41422
rect 90302 41346 90354 41358
rect 53342 41298 53394 41310
rect 53342 41234 53394 41246
rect 53790 41298 53842 41310
rect 53790 41234 53842 41246
rect 54238 41298 54290 41310
rect 54238 41234 54290 41246
rect 55134 41298 55186 41310
rect 55134 41234 55186 41246
rect 56590 41298 56642 41310
rect 56590 41234 56642 41246
rect 56926 41298 56978 41310
rect 65550 41298 65602 41310
rect 62178 41246 62190 41298
rect 62242 41246 62254 41298
rect 64306 41246 64318 41298
rect 64370 41246 64382 41298
rect 56926 41234 56978 41246
rect 65550 41234 65602 41246
rect 68686 41298 68738 41310
rect 70366 41298 70418 41310
rect 69458 41246 69470 41298
rect 69522 41246 69534 41298
rect 68686 41234 68738 41246
rect 70366 41234 70418 41246
rect 70814 41298 70866 41310
rect 70814 41234 70866 41246
rect 72270 41298 72322 41310
rect 72270 41234 72322 41246
rect 72718 41298 72770 41310
rect 72718 41234 72770 41246
rect 75854 41298 75906 41310
rect 75854 41234 75906 41246
rect 84254 41298 84306 41310
rect 86706 41246 86718 41298
rect 86770 41246 86782 41298
rect 93202 41246 93214 41298
rect 93266 41246 93278 41298
rect 95330 41246 95342 41298
rect 95394 41246 95406 41298
rect 84254 41234 84306 41246
rect 50766 41186 50818 41198
rect 58606 41186 58658 41198
rect 60286 41186 60338 41198
rect 65998 41186 66050 41198
rect 52546 41134 52558 41186
rect 52610 41134 52622 41186
rect 57698 41134 57710 41186
rect 57762 41134 57774 41186
rect 59714 41134 59726 41186
rect 59778 41134 59790 41186
rect 64978 41134 64990 41186
rect 65042 41134 65054 41186
rect 50766 41122 50818 41134
rect 58606 41122 58658 41134
rect 60286 41122 60338 41134
rect 65998 41122 66050 41134
rect 67678 41186 67730 41198
rect 73838 41186 73890 41198
rect 82462 41186 82514 41198
rect 90638 41186 90690 41198
rect 97134 41186 97186 41198
rect 71810 41134 71822 41186
rect 71874 41134 71886 41186
rect 77522 41134 77534 41186
rect 77586 41134 77598 41186
rect 85810 41134 85822 41186
rect 85874 41134 85886 41186
rect 89618 41134 89630 41186
rect 89682 41134 89694 41186
rect 91298 41134 91310 41186
rect 91362 41134 91374 41186
rect 96114 41134 96126 41186
rect 96178 41134 96190 41186
rect 97570 41134 97582 41186
rect 97634 41134 97646 41186
rect 67678 41122 67730 41134
rect 73838 41122 73890 41134
rect 82462 41122 82514 41134
rect 90638 41122 90690 41134
rect 97134 41122 97186 41134
rect 49534 41074 49586 41086
rect 49534 41010 49586 41022
rect 49870 41074 49922 41086
rect 49870 41010 49922 41022
rect 50430 41074 50482 41086
rect 50430 41010 50482 41022
rect 51438 41074 51490 41086
rect 54686 41074 54738 41086
rect 52322 41022 52334 41074
rect 52386 41022 52398 41074
rect 51438 41010 51490 41022
rect 54686 41010 54738 41022
rect 57934 41074 57986 41086
rect 67342 41074 67394 41086
rect 77310 41074 77362 41086
rect 59490 41022 59502 41074
rect 59554 41022 59566 41074
rect 74050 41022 74062 41074
rect 74114 41022 74126 41074
rect 74610 41022 74622 41074
rect 74674 41022 74686 41074
rect 57934 41010 57986 41022
rect 67342 41010 67394 41022
rect 77310 41010 77362 41022
rect 78990 41074 79042 41086
rect 78990 41010 79042 41022
rect 81566 41074 81618 41086
rect 85598 41074 85650 41086
rect 92430 41074 92482 41086
rect 82674 41022 82686 41074
rect 82738 41022 82750 41074
rect 83234 41022 83246 41074
rect 83298 41022 83310 41074
rect 88834 41022 88846 41074
rect 88898 41022 88910 41074
rect 91186 41022 91198 41074
rect 91250 41022 91262 41074
rect 81566 41010 81618 41022
rect 85598 41010 85650 41022
rect 92430 41010 92482 41022
rect 96798 41074 96850 41086
rect 97906 41022 97918 41074
rect 97970 41022 97982 41074
rect 96798 41010 96850 41022
rect 69918 40962 69970 40974
rect 69918 40898 69970 40910
rect 73502 40962 73554 40974
rect 73502 40898 73554 40910
rect 75294 40962 75346 40974
rect 75294 40898 75346 40910
rect 76302 40962 76354 40974
rect 76302 40898 76354 40910
rect 79326 40962 79378 40974
rect 79326 40898 79378 40910
rect 83806 40962 83858 40974
rect 83806 40898 83858 40910
rect 92094 40962 92146 40974
rect 92094 40898 92146 40910
rect 1344 40794 98560 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 98560 40794
rect 1344 40708 98560 40742
rect 62190 40626 62242 40638
rect 62190 40562 62242 40574
rect 62750 40626 62802 40638
rect 62750 40562 62802 40574
rect 64542 40626 64594 40638
rect 64542 40562 64594 40574
rect 70702 40626 70754 40638
rect 70702 40562 70754 40574
rect 71262 40626 71314 40638
rect 71262 40562 71314 40574
rect 72270 40626 72322 40638
rect 72270 40562 72322 40574
rect 74174 40626 74226 40638
rect 74174 40562 74226 40574
rect 74622 40626 74674 40638
rect 74622 40562 74674 40574
rect 89294 40626 89346 40638
rect 89294 40562 89346 40574
rect 98030 40626 98082 40638
rect 98030 40562 98082 40574
rect 73390 40514 73442 40526
rect 96126 40514 96178 40526
rect 53330 40462 53342 40514
rect 53394 40462 53406 40514
rect 59602 40462 59614 40514
rect 59666 40462 59678 40514
rect 63522 40462 63534 40514
rect 63586 40462 63598 40514
rect 63970 40462 63982 40514
rect 64034 40462 64046 40514
rect 88162 40462 88174 40514
rect 88226 40462 88238 40514
rect 73390 40450 73442 40462
rect 96126 40450 96178 40462
rect 97246 40514 97298 40526
rect 97246 40450 97298 40462
rect 56030 40402 56082 40414
rect 55570 40350 55582 40402
rect 55634 40350 55646 40402
rect 56030 40338 56082 40350
rect 58158 40402 58210 40414
rect 65326 40402 65378 40414
rect 81230 40402 81282 40414
rect 58930 40350 58942 40402
rect 58994 40350 59006 40402
rect 67442 40350 67454 40402
rect 67506 40350 67518 40402
rect 73602 40350 73614 40402
rect 73666 40350 73678 40402
rect 80434 40350 80446 40402
rect 80498 40350 80510 40402
rect 58158 40338 58210 40350
rect 65326 40338 65378 40350
rect 81230 40338 81282 40350
rect 82686 40402 82738 40414
rect 83906 40350 83918 40402
rect 83970 40350 83982 40402
rect 89506 40350 89518 40402
rect 89570 40350 89582 40402
rect 95666 40350 95678 40402
rect 95730 40350 95742 40402
rect 97458 40350 97470 40402
rect 97522 40350 97534 40402
rect 82686 40338 82738 40350
rect 64206 40290 64258 40302
rect 61730 40238 61742 40290
rect 61794 40238 61806 40290
rect 68114 40238 68126 40290
rect 68178 40238 68190 40290
rect 70242 40238 70254 40290
rect 70306 40238 70318 40290
rect 71698 40238 71710 40290
rect 71762 40238 71774 40290
rect 77746 40238 77758 40290
rect 77810 40238 77822 40290
rect 90850 40238 90862 40290
rect 90914 40238 90926 40290
rect 64206 40226 64258 40238
rect 1344 40010 98560 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 98560 40010
rect 1344 39924 98560 39958
rect 70702 39730 70754 39742
rect 77198 39730 77250 39742
rect 85150 39730 85202 39742
rect 93326 39730 93378 39742
rect 64978 39678 64990 39730
rect 65042 39678 65054 39730
rect 72706 39678 72718 39730
rect 72770 39678 72782 39730
rect 74834 39678 74846 39730
rect 74898 39678 74910 39730
rect 75842 39678 75854 39730
rect 75906 39678 75918 39730
rect 79202 39678 79214 39730
rect 79266 39678 79278 39730
rect 81330 39678 81342 39730
rect 81394 39678 81406 39730
rect 87938 39678 87950 39730
rect 88002 39678 88014 39730
rect 94882 39678 94894 39730
rect 94946 39678 94958 39730
rect 97010 39678 97022 39730
rect 97074 39678 97086 39730
rect 70702 39666 70754 39678
rect 77198 39666 77250 39678
rect 85150 39666 85202 39678
rect 93326 39666 93378 39678
rect 53454 39618 53506 39630
rect 53454 39554 53506 39566
rect 61742 39618 61794 39630
rect 69694 39618 69746 39630
rect 62290 39566 62302 39618
rect 62354 39566 62366 39618
rect 61742 39554 61794 39566
rect 69694 39554 69746 39566
rect 70254 39618 70306 39630
rect 75406 39618 75458 39630
rect 72034 39566 72046 39618
rect 72098 39566 72110 39618
rect 70254 39554 70306 39566
rect 75406 39554 75458 39566
rect 76414 39618 76466 39630
rect 83246 39618 83298 39630
rect 78418 39566 78430 39618
rect 78482 39566 78494 39618
rect 82338 39566 82350 39618
rect 82402 39566 82414 39618
rect 76414 39554 76466 39566
rect 83246 39554 83298 39566
rect 83582 39618 83634 39630
rect 93886 39618 93938 39630
rect 84130 39566 84142 39618
rect 84194 39566 84206 39618
rect 90850 39566 90862 39618
rect 90914 39566 90926 39618
rect 97794 39566 97806 39618
rect 97858 39566 97870 39618
rect 83582 39554 83634 39566
rect 93886 39554 93938 39566
rect 51102 39506 51154 39518
rect 51102 39442 51154 39454
rect 51438 39506 51490 39518
rect 51438 39442 51490 39454
rect 55806 39506 55858 39518
rect 55806 39442 55858 39454
rect 59950 39506 60002 39518
rect 59950 39442 60002 39454
rect 68238 39506 68290 39518
rect 68238 39442 68290 39454
rect 68574 39506 68626 39518
rect 84354 39454 84366 39506
rect 84418 39454 84430 39506
rect 90066 39454 90078 39506
rect 90130 39454 90142 39506
rect 68574 39442 68626 39454
rect 50542 39394 50594 39406
rect 50542 39330 50594 39342
rect 55470 39394 55522 39406
rect 55470 39330 55522 39342
rect 59614 39394 59666 39406
rect 59614 39330 59666 39342
rect 61294 39394 61346 39406
rect 61294 39330 61346 39342
rect 77870 39394 77922 39406
rect 77870 39330 77922 39342
rect 82574 39394 82626 39406
rect 82574 39330 82626 39342
rect 94222 39394 94274 39406
rect 94222 39330 94274 39342
rect 1344 39226 98560 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 98560 39226
rect 1344 39140 98560 39174
rect 62190 39058 62242 39070
rect 62190 38994 62242 39006
rect 69694 39058 69746 39070
rect 69694 38994 69746 39006
rect 71374 39058 71426 39070
rect 71374 38994 71426 39006
rect 78990 39058 79042 39070
rect 78990 38994 79042 39006
rect 81342 39058 81394 39070
rect 81342 38994 81394 39006
rect 85822 39058 85874 39070
rect 85822 38994 85874 39006
rect 88510 39058 88562 39070
rect 88510 38994 88562 39006
rect 89630 39058 89682 39070
rect 89630 38994 89682 39006
rect 94558 39058 94610 39070
rect 94558 38994 94610 39006
rect 96350 39058 96402 39070
rect 96350 38994 96402 39006
rect 97134 39058 97186 39070
rect 97134 38994 97186 39006
rect 97582 39058 97634 39070
rect 97582 38994 97634 39006
rect 50318 38946 50370 38958
rect 53006 38946 53058 38958
rect 63982 38946 64034 38958
rect 74846 38946 74898 38958
rect 90526 38946 90578 38958
rect 52210 38894 52222 38946
rect 52274 38894 52286 38946
rect 54562 38894 54574 38946
rect 54626 38894 54638 38946
rect 59378 38894 59390 38946
rect 59442 38894 59454 38946
rect 63074 38894 63086 38946
rect 63138 38894 63150 38946
rect 70802 38894 70814 38946
rect 70866 38894 70878 38946
rect 76178 38894 76190 38946
rect 76242 38894 76254 38946
rect 80098 38894 80110 38946
rect 80162 38894 80174 38946
rect 83234 38894 83246 38946
rect 83298 38894 83310 38946
rect 91858 38894 91870 38946
rect 91922 38894 91934 38946
rect 95442 38894 95454 38946
rect 95506 38894 95518 38946
rect 50318 38882 50370 38894
rect 53006 38882 53058 38894
rect 63982 38882 64034 38894
rect 74846 38882 74898 38894
rect 90526 38882 90578 38894
rect 50654 38834 50706 38846
rect 50654 38770 50706 38782
rect 51326 38834 51378 38846
rect 62526 38834 62578 38846
rect 70030 38834 70082 38846
rect 90190 38834 90242 38846
rect 96014 38834 96066 38846
rect 52434 38782 52446 38834
rect 52498 38782 52510 38834
rect 53778 38782 53790 38834
rect 53842 38782 53854 38834
rect 58706 38782 58718 38834
rect 58770 38782 58782 38834
rect 63186 38782 63198 38834
rect 63250 38782 63262 38834
rect 64194 38782 64206 38834
rect 64258 38782 64270 38834
rect 65538 38782 65550 38834
rect 65602 38782 65614 38834
rect 70690 38782 70702 38834
rect 70754 38782 70766 38834
rect 74610 38782 74622 38834
rect 74674 38782 74686 38834
rect 75506 38782 75518 38834
rect 75570 38782 75582 38834
rect 79986 38782 79998 38834
rect 80050 38782 80062 38834
rect 82562 38782 82574 38834
rect 82626 38782 82638 38834
rect 89394 38782 89406 38834
rect 89458 38782 89470 38834
rect 91186 38782 91198 38834
rect 91250 38782 91262 38834
rect 95218 38782 95230 38834
rect 95282 38782 95294 38834
rect 51326 38770 51378 38782
rect 62526 38770 62578 38782
rect 70030 38770 70082 38782
rect 90190 38770 90242 38782
rect 96014 38770 96066 38782
rect 71822 38722 71874 38734
rect 79326 38722 79378 38734
rect 98030 38722 98082 38734
rect 56690 38670 56702 38722
rect 56754 38670 56766 38722
rect 61506 38670 61518 38722
rect 61570 38670 61582 38722
rect 66210 38670 66222 38722
rect 66274 38670 66286 38722
rect 68338 38670 68350 38722
rect 68402 38670 68414 38722
rect 78306 38670 78318 38722
rect 78370 38670 78382 38722
rect 85362 38670 85374 38722
rect 85426 38670 85438 38722
rect 93986 38670 93998 38722
rect 94050 38670 94062 38722
rect 71822 38658 71874 38670
rect 79326 38658 79378 38670
rect 98030 38658 98082 38670
rect 51662 38610 51714 38622
rect 51662 38546 51714 38558
rect 1344 38442 98560 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 98560 38442
rect 1344 38356 98560 38390
rect 56366 38274 56418 38286
rect 56366 38210 56418 38222
rect 56702 38274 56754 38286
rect 56702 38210 56754 38222
rect 74846 38274 74898 38286
rect 74846 38210 74898 38222
rect 75182 38274 75234 38286
rect 75182 38210 75234 38222
rect 53454 38162 53506 38174
rect 50530 38110 50542 38162
rect 50594 38110 50606 38162
rect 52658 38110 52670 38162
rect 52722 38110 52734 38162
rect 53454 38098 53506 38110
rect 53790 38162 53842 38174
rect 53790 38098 53842 38110
rect 61518 38162 61570 38174
rect 65550 38162 65602 38174
rect 62850 38110 62862 38162
rect 62914 38110 62926 38162
rect 64978 38110 64990 38162
rect 65042 38110 65054 38162
rect 61518 38098 61570 38110
rect 65550 38098 65602 38110
rect 69246 38162 69298 38174
rect 69246 38098 69298 38110
rect 69694 38162 69746 38174
rect 69694 38098 69746 38110
rect 76526 38162 76578 38174
rect 76526 38098 76578 38110
rect 78990 38162 79042 38174
rect 85150 38162 85202 38174
rect 84242 38110 84254 38162
rect 84306 38110 84318 38162
rect 78990 38098 79042 38110
rect 85150 38098 85202 38110
rect 93326 38162 93378 38174
rect 98030 38162 98082 38174
rect 97570 38110 97582 38162
rect 97634 38110 97646 38162
rect 93326 38098 93378 38110
rect 98030 38098 98082 38110
rect 67566 38050 67618 38062
rect 77310 38050 77362 38062
rect 48962 37998 48974 38050
rect 49026 37998 49038 38050
rect 49746 37998 49758 38050
rect 49810 37998 49822 38050
rect 57362 37998 57374 38050
rect 57426 37998 57438 38050
rect 62178 37998 62190 38050
rect 62242 37998 62254 38050
rect 68338 37998 68350 38050
rect 68402 37998 68414 38050
rect 75842 37998 75854 38050
rect 75906 37998 75918 38050
rect 67566 37986 67618 37998
rect 77310 37986 77362 37998
rect 77870 38050 77922 38062
rect 77870 37986 77922 37998
rect 78542 38050 78594 38062
rect 91646 38050 91698 38062
rect 81442 37998 81454 38050
rect 81506 37998 81518 38050
rect 89170 37998 89182 38050
rect 89234 37998 89246 38050
rect 90962 37998 90974 38050
rect 91026 37998 91038 38050
rect 94658 37998 94670 38050
rect 94722 37998 94734 38050
rect 78542 37986 78594 37998
rect 91646 37986 91698 37998
rect 1822 37938 1874 37950
rect 1822 37874 1874 37886
rect 2158 37938 2210 37950
rect 66222 37938 66274 37950
rect 57250 37886 57262 37938
rect 57314 37886 57326 37938
rect 2158 37874 2210 37886
rect 66222 37874 66274 37886
rect 66558 37938 66610 37950
rect 66558 37874 66610 37886
rect 67230 37938 67282 37950
rect 93774 37938 93826 37950
rect 68226 37886 68238 37938
rect 68290 37886 68302 37938
rect 75954 37886 75966 37938
rect 76018 37886 76030 37938
rect 82114 37886 82126 37938
rect 82178 37886 82190 37938
rect 90850 37886 90862 37938
rect 90914 37886 90926 37938
rect 67230 37874 67282 37886
rect 93774 37874 93826 37886
rect 94110 37938 94162 37950
rect 95442 37886 95454 37938
rect 95506 37886 95518 37938
rect 94110 37874 94162 37886
rect 49198 37826 49250 37838
rect 49198 37762 49250 37774
rect 55694 37826 55746 37838
rect 55694 37762 55746 37774
rect 58046 37826 58098 37838
rect 58046 37762 58098 37774
rect 88510 37826 88562 37838
rect 88510 37762 88562 37774
rect 89406 37826 89458 37838
rect 89406 37762 89458 37774
rect 89854 37826 89906 37838
rect 89854 37762 89906 37774
rect 91982 37826 92034 37838
rect 91982 37762 92034 37774
rect 1344 37658 98560 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 98560 37658
rect 1344 37572 98560 37606
rect 1822 37490 1874 37502
rect 1822 37426 1874 37438
rect 52894 37490 52946 37502
rect 52894 37426 52946 37438
rect 59390 37490 59442 37502
rect 59390 37426 59442 37438
rect 59838 37490 59890 37502
rect 59838 37426 59890 37438
rect 63422 37490 63474 37502
rect 63422 37426 63474 37438
rect 65326 37490 65378 37502
rect 65326 37426 65378 37438
rect 65774 37490 65826 37502
rect 65774 37426 65826 37438
rect 74174 37490 74226 37502
rect 74174 37426 74226 37438
rect 75294 37490 75346 37502
rect 75294 37426 75346 37438
rect 77086 37490 77138 37502
rect 77086 37426 77138 37438
rect 81902 37490 81954 37502
rect 81902 37426 81954 37438
rect 93886 37490 93938 37502
rect 93886 37426 93938 37438
rect 94222 37490 94274 37502
rect 94222 37426 94274 37438
rect 96350 37490 96402 37502
rect 96350 37426 96402 37438
rect 56702 37378 56754 37390
rect 77870 37378 77922 37390
rect 92766 37378 92818 37390
rect 50306 37326 50318 37378
rect 50370 37326 50382 37378
rect 58818 37326 58830 37378
rect 58882 37326 58894 37378
rect 64306 37326 64318 37378
rect 64370 37326 64382 37378
rect 75842 37326 75854 37378
rect 75906 37326 75918 37378
rect 76402 37326 76414 37378
rect 76466 37326 76478 37378
rect 83794 37326 83806 37378
rect 83858 37326 83870 37378
rect 91410 37326 91422 37378
rect 91474 37326 91486 37378
rect 56702 37314 56754 37326
rect 77870 37314 77922 37326
rect 92766 37314 92818 37326
rect 93102 37378 93154 37390
rect 95330 37326 95342 37378
rect 95394 37326 95406 37378
rect 93102 37314 93154 37326
rect 57710 37266 57762 37278
rect 75630 37266 75682 37278
rect 49634 37214 49646 37266
rect 49698 37214 49710 37266
rect 56466 37214 56478 37266
rect 56530 37214 56542 37266
rect 58706 37214 58718 37266
rect 58770 37214 58782 37266
rect 64418 37214 64430 37266
rect 64482 37214 64494 37266
rect 66770 37214 66782 37266
rect 66834 37214 66846 37266
rect 57710 37202 57762 37214
rect 75630 37202 75682 37214
rect 82238 37266 82290 37278
rect 82238 37202 82290 37214
rect 82910 37266 82962 37278
rect 82910 37202 82962 37214
rect 83246 37266 83298 37278
rect 96014 37266 96066 37278
rect 83906 37214 83918 37266
rect 83970 37214 83982 37266
rect 92194 37214 92206 37266
rect 92258 37214 92270 37266
rect 95442 37214 95454 37266
rect 95506 37214 95518 37266
rect 83246 37202 83298 37214
rect 96014 37202 96066 37214
rect 70142 37154 70194 37166
rect 52434 37102 52446 37154
rect 52498 37102 52510 37154
rect 67442 37102 67454 37154
rect 67506 37102 67518 37154
rect 69570 37102 69582 37154
rect 69634 37102 69646 37154
rect 70142 37090 70194 37102
rect 74622 37154 74674 37166
rect 74622 37090 74674 37102
rect 77422 37154 77474 37166
rect 77422 37090 77474 37102
rect 84590 37154 84642 37166
rect 97134 37154 97186 37166
rect 89282 37102 89294 37154
rect 89346 37102 89358 37154
rect 84590 37090 84642 37102
rect 97134 37090 97186 37102
rect 58046 37042 58098 37054
rect 58046 36978 58098 36990
rect 63758 37042 63810 37054
rect 63758 36978 63810 36990
rect 1344 36874 98560 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 98560 36874
rect 1344 36788 98560 36822
rect 51102 36706 51154 36718
rect 51102 36642 51154 36654
rect 51438 36706 51490 36718
rect 69806 36706 69858 36718
rect 64866 36654 64878 36706
rect 64930 36703 64942 36706
rect 65426 36703 65438 36706
rect 64930 36657 65438 36703
rect 64930 36654 64942 36657
rect 65426 36654 65438 36657
rect 65490 36654 65502 36706
rect 51438 36642 51490 36654
rect 69806 36642 69858 36654
rect 95230 36706 95282 36718
rect 95230 36642 95282 36654
rect 95566 36706 95618 36718
rect 95566 36642 95618 36654
rect 53790 36594 53842 36606
rect 61518 36594 61570 36606
rect 56802 36542 56814 36594
rect 56866 36542 56878 36594
rect 58930 36542 58942 36594
rect 58994 36542 59006 36594
rect 53790 36530 53842 36542
rect 61518 36530 61570 36542
rect 64990 36594 65042 36606
rect 64990 36530 65042 36542
rect 65438 36594 65490 36606
rect 65438 36530 65490 36542
rect 71150 36594 71202 36606
rect 71150 36530 71202 36542
rect 73390 36594 73442 36606
rect 77198 36594 77250 36606
rect 74274 36542 74286 36594
rect 74338 36542 74350 36594
rect 73390 36530 73442 36542
rect 77198 36530 77250 36542
rect 77646 36594 77698 36606
rect 77646 36530 77698 36542
rect 82574 36594 82626 36606
rect 82574 36530 82626 36542
rect 87054 36594 87106 36606
rect 93214 36594 93266 36606
rect 89506 36542 89518 36594
rect 89570 36542 89582 36594
rect 91634 36542 91646 36594
rect 91698 36542 91710 36594
rect 87054 36530 87106 36542
rect 93214 36530 93266 36542
rect 96910 36594 96962 36606
rect 96910 36530 96962 36542
rect 53342 36482 53394 36494
rect 73838 36482 73890 36494
rect 52210 36430 52222 36482
rect 52274 36430 52286 36482
rect 56130 36430 56142 36482
rect 56194 36430 56206 36482
rect 70578 36430 70590 36482
rect 70642 36430 70654 36482
rect 53342 36418 53394 36430
rect 73838 36418 73890 36430
rect 74958 36482 75010 36494
rect 76078 36482 76130 36494
rect 93774 36482 93826 36494
rect 75394 36430 75406 36482
rect 75458 36430 75470 36482
rect 92418 36430 92430 36482
rect 92482 36430 92494 36482
rect 94322 36430 94334 36482
rect 94386 36430 94398 36482
rect 74958 36418 75010 36430
rect 76078 36418 76130 36430
rect 93774 36418 93826 36430
rect 59502 36370 59554 36382
rect 52098 36318 52110 36370
rect 52162 36318 52174 36370
rect 59502 36306 59554 36318
rect 68014 36370 68066 36382
rect 68014 36306 68066 36318
rect 68350 36370 68402 36382
rect 68350 36306 68402 36318
rect 69470 36370 69522 36382
rect 71598 36370 71650 36382
rect 70354 36318 70366 36370
rect 70418 36318 70430 36370
rect 69470 36306 69522 36318
rect 71598 36306 71650 36318
rect 76414 36370 76466 36382
rect 95778 36318 95790 36370
rect 95842 36318 95854 36370
rect 96226 36318 96238 36370
rect 96290 36318 96302 36370
rect 76414 36306 76466 36318
rect 54238 36258 54290 36270
rect 54238 36194 54290 36206
rect 59838 36258 59890 36270
rect 59838 36194 59890 36206
rect 60286 36258 60338 36270
rect 60286 36194 60338 36206
rect 94558 36258 94610 36270
rect 94558 36194 94610 36206
rect 1344 36090 98560 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 98560 36090
rect 1344 36004 98560 36038
rect 55246 35922 55298 35934
rect 55246 35858 55298 35870
rect 56702 35922 56754 35934
rect 56702 35858 56754 35870
rect 59054 35922 59106 35934
rect 59054 35858 59106 35870
rect 59726 35922 59778 35934
rect 59726 35858 59778 35870
rect 61070 35922 61122 35934
rect 61070 35858 61122 35870
rect 64542 35922 64594 35934
rect 64542 35858 64594 35870
rect 74062 35922 74114 35934
rect 74062 35858 74114 35870
rect 77310 35922 77362 35934
rect 77310 35858 77362 35870
rect 81230 35922 81282 35934
rect 81230 35858 81282 35870
rect 81678 35922 81730 35934
rect 81678 35858 81730 35870
rect 82462 35922 82514 35934
rect 82462 35858 82514 35870
rect 84478 35922 84530 35934
rect 84478 35858 84530 35870
rect 84926 35922 84978 35934
rect 84926 35858 84978 35870
rect 89406 35922 89458 35934
rect 89406 35858 89458 35870
rect 60622 35810 60674 35822
rect 71710 35810 71762 35822
rect 76526 35810 76578 35822
rect 54114 35758 54126 35810
rect 54178 35758 54190 35810
rect 54450 35758 54462 35810
rect 54514 35758 54526 35810
rect 58034 35758 58046 35810
rect 58098 35758 58110 35810
rect 58482 35758 58494 35810
rect 58546 35758 58558 35810
rect 61954 35758 61966 35810
rect 62018 35758 62030 35810
rect 62514 35758 62526 35810
rect 62578 35758 62590 35810
rect 74946 35758 74958 35810
rect 75010 35758 75022 35810
rect 60622 35746 60674 35758
rect 71710 35746 71762 35758
rect 76526 35746 76578 35758
rect 83358 35810 83410 35822
rect 87614 35810 87666 35822
rect 86146 35758 86158 35810
rect 86210 35758 86222 35810
rect 86706 35758 86718 35810
rect 86770 35758 86782 35810
rect 83358 35746 83410 35758
rect 87614 35746 87666 35758
rect 88510 35810 88562 35822
rect 97134 35810 97186 35822
rect 89954 35758 89966 35810
rect 90018 35758 90030 35810
rect 90290 35758 90302 35810
rect 90354 35758 90366 35810
rect 88510 35746 88562 35758
rect 97134 35746 97186 35758
rect 60286 35698 60338 35710
rect 49970 35646 49982 35698
rect 50034 35646 50046 35698
rect 60286 35634 60338 35646
rect 62750 35698 62802 35710
rect 62750 35634 62802 35646
rect 63086 35698 63138 35710
rect 89742 35698 89794 35710
rect 71922 35646 71934 35698
rect 71986 35646 71998 35698
rect 74722 35646 74734 35698
rect 74786 35646 74798 35698
rect 76738 35646 76750 35698
rect 76802 35646 76814 35698
rect 83122 35646 83134 35698
rect 83186 35646 83198 35698
rect 87826 35646 87838 35698
rect 87890 35646 87902 35698
rect 96450 35646 96462 35698
rect 96514 35646 96526 35698
rect 63086 35634 63138 35646
rect 89742 35634 89794 35646
rect 63646 35586 63698 35598
rect 50754 35534 50766 35586
rect 50818 35534 50830 35586
rect 52882 35534 52894 35586
rect 52946 35534 52958 35586
rect 63646 35522 63698 35534
rect 66670 35586 66722 35598
rect 66670 35522 66722 35534
rect 72606 35586 72658 35598
rect 72606 35522 72658 35534
rect 73502 35586 73554 35598
rect 73502 35522 73554 35534
rect 75854 35586 75906 35598
rect 94434 35534 94446 35586
rect 94498 35534 94510 35586
rect 75854 35522 75906 35534
rect 53566 35474 53618 35486
rect 53566 35410 53618 35422
rect 53902 35474 53954 35486
rect 53902 35410 53954 35422
rect 58718 35474 58770 35486
rect 58718 35410 58770 35422
rect 75518 35474 75570 35486
rect 85598 35474 85650 35486
rect 84466 35422 84478 35474
rect 84530 35471 84542 35474
rect 85250 35471 85262 35474
rect 84530 35425 85262 35471
rect 84530 35422 84542 35425
rect 85250 35422 85262 35425
rect 85314 35422 85326 35474
rect 75518 35410 75570 35422
rect 85598 35410 85650 35422
rect 85934 35474 85986 35486
rect 85934 35410 85986 35422
rect 1344 35306 98560 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 98560 35306
rect 1344 35220 98560 35254
rect 71822 35138 71874 35150
rect 71822 35074 71874 35086
rect 53454 35026 53506 35038
rect 66670 35026 66722 35038
rect 88622 35026 88674 35038
rect 52658 34974 52670 35026
rect 52722 34974 52734 35026
rect 57362 34974 57374 35026
rect 57426 34974 57438 35026
rect 62178 34974 62190 35026
rect 62242 34974 62254 35026
rect 64306 34974 64318 35026
rect 64370 34974 64382 35026
rect 74386 34974 74398 35026
rect 74450 34974 74462 35026
rect 76514 34974 76526 35026
rect 76578 34974 76590 35026
rect 81666 34974 81678 35026
rect 81730 34974 81742 35026
rect 88162 34974 88174 35026
rect 88226 34974 88238 35026
rect 53454 34962 53506 34974
rect 66670 34962 66722 34974
rect 88622 34962 88674 34974
rect 90302 35026 90354 35038
rect 97234 34974 97246 35026
rect 97298 34974 97310 35026
rect 90302 34962 90354 34974
rect 65326 34914 65378 34926
rect 67678 34914 67730 34926
rect 69694 34914 69746 34926
rect 49858 34862 49870 34914
rect 49922 34862 49934 34914
rect 56802 34862 56814 34914
rect 56866 34862 56878 34914
rect 61394 34862 61406 34914
rect 61458 34862 61470 34914
rect 66098 34862 66110 34914
rect 66162 34862 66174 34914
rect 68450 34862 68462 34914
rect 68514 34862 68526 34914
rect 65326 34850 65378 34862
rect 67678 34850 67730 34862
rect 69694 34850 69746 34862
rect 72158 34914 72210 34926
rect 77310 34914 77362 34926
rect 82686 34914 82738 34926
rect 91646 34914 91698 34926
rect 73714 34862 73726 34914
rect 73778 34862 73790 34914
rect 78754 34862 78766 34914
rect 78818 34862 78830 34914
rect 84242 34862 84254 34914
rect 84306 34862 84318 34914
rect 85250 34862 85262 34914
rect 85314 34862 85326 34914
rect 90962 34862 90974 34914
rect 91026 34862 91038 34914
rect 94434 34862 94446 34914
rect 94498 34862 94510 34914
rect 72158 34850 72210 34862
rect 77310 34850 77362 34862
rect 82686 34850 82738 34862
rect 91646 34850 91698 34862
rect 54350 34802 54402 34814
rect 50530 34750 50542 34802
rect 50594 34750 50606 34802
rect 54350 34738 54402 34750
rect 54686 34802 54738 34814
rect 71150 34802 71202 34814
rect 84478 34802 84530 34814
rect 65874 34750 65886 34802
rect 65938 34750 65950 34802
rect 68226 34750 68238 34802
rect 68290 34750 68302 34802
rect 72370 34750 72382 34802
rect 72434 34750 72446 34802
rect 72706 34750 72718 34802
rect 72770 34750 72782 34802
rect 79538 34750 79550 34802
rect 79602 34750 79614 34802
rect 82898 34750 82910 34802
rect 82962 34750 82974 34802
rect 83234 34750 83246 34802
rect 83298 34750 83310 34802
rect 86034 34750 86046 34802
rect 86098 34750 86110 34802
rect 90850 34750 90862 34802
rect 90914 34750 90926 34802
rect 95106 34750 95118 34802
rect 95170 34750 95182 34802
rect 54686 34738 54738 34750
rect 71150 34738 71202 34750
rect 84478 34738 84530 34750
rect 53790 34690 53842 34702
rect 53790 34626 53842 34638
rect 64990 34690 65042 34702
rect 64990 34626 65042 34638
rect 67342 34690 67394 34702
rect 67342 34626 67394 34638
rect 69358 34690 69410 34702
rect 69358 34626 69410 34638
rect 70814 34690 70866 34702
rect 70814 34626 70866 34638
rect 82350 34690 82402 34702
rect 82350 34626 82402 34638
rect 89854 34690 89906 34702
rect 89854 34626 89906 34638
rect 91982 34690 92034 34702
rect 91982 34626 92034 34638
rect 1344 34522 98560 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 98560 34522
rect 1344 34436 98560 34470
rect 50990 34354 51042 34366
rect 50990 34290 51042 34302
rect 64542 34354 64594 34366
rect 64542 34290 64594 34302
rect 66222 34354 66274 34366
rect 66222 34290 66274 34302
rect 73502 34354 73554 34366
rect 73502 34290 73554 34302
rect 75294 34354 75346 34366
rect 75294 34290 75346 34302
rect 79550 34354 79602 34366
rect 79550 34290 79602 34302
rect 93662 34354 93714 34366
rect 93662 34290 93714 34302
rect 94558 34354 94610 34366
rect 94558 34290 94610 34302
rect 95230 34354 95282 34366
rect 95230 34290 95282 34302
rect 97134 34354 97186 34366
rect 97134 34290 97186 34302
rect 51326 34242 51378 34254
rect 65438 34242 65490 34254
rect 52994 34190 53006 34242
rect 53058 34190 53070 34242
rect 59602 34190 59614 34242
rect 59666 34190 59678 34242
rect 51326 34178 51378 34190
rect 65438 34178 65490 34190
rect 65774 34242 65826 34254
rect 79886 34242 79938 34254
rect 92766 34242 92818 34254
rect 70130 34190 70142 34242
rect 70194 34190 70206 34242
rect 74386 34190 74398 34242
rect 74450 34190 74462 34242
rect 87938 34190 87950 34242
rect 88002 34190 88014 34242
rect 88162 34190 88174 34242
rect 88226 34190 88238 34242
rect 65774 34178 65826 34190
rect 79886 34178 79938 34190
rect 92766 34178 92818 34190
rect 93102 34242 93154 34254
rect 95778 34190 95790 34242
rect 95842 34190 95854 34242
rect 96114 34190 96126 34242
rect 96178 34190 96190 34242
rect 93102 34178 93154 34190
rect 52334 34130 52386 34142
rect 73838 34130 73890 34142
rect 95566 34130 95618 34142
rect 53106 34078 53118 34130
rect 53170 34078 53182 34130
rect 53890 34078 53902 34130
rect 53954 34078 53966 34130
rect 60274 34078 60286 34130
rect 60338 34078 60350 34130
rect 60946 34078 60958 34130
rect 61010 34078 61022 34130
rect 67218 34078 67230 34130
rect 67282 34078 67294 34130
rect 74610 34078 74622 34130
rect 74674 34078 74686 34130
rect 78754 34078 78766 34130
rect 78818 34078 78830 34130
rect 86594 34078 86606 34130
rect 86658 34078 86670 34130
rect 89394 34078 89406 34130
rect 89458 34078 89470 34130
rect 94322 34078 94334 34130
rect 94386 34078 94398 34130
rect 52334 34066 52386 34078
rect 73838 34066 73890 34078
rect 95566 34066 95618 34078
rect 87614 34018 87666 34030
rect 54562 33966 54574 34018
rect 54626 33966 54638 34018
rect 56690 33966 56702 34018
rect 56754 33966 56766 34018
rect 57474 33966 57486 34018
rect 57538 33966 57550 34018
rect 61730 33966 61742 34018
rect 61794 33966 61806 34018
rect 63858 33966 63870 34018
rect 63922 33966 63934 34018
rect 75954 33966 75966 34018
rect 76018 33966 76030 34018
rect 78082 33966 78094 34018
rect 78146 33966 78158 34018
rect 82450 33966 82462 34018
rect 82514 33966 82526 34018
rect 90066 33966 90078 34018
rect 90130 33966 90142 34018
rect 92194 33966 92206 34018
rect 92258 33966 92270 34018
rect 87614 33954 87666 33966
rect 51998 33906 52050 33918
rect 51998 33842 52050 33854
rect 87278 33906 87330 33918
rect 87278 33842 87330 33854
rect 1344 33738 98560 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 98560 33738
rect 1344 33652 98560 33686
rect 82126 33570 82178 33582
rect 72818 33518 72830 33570
rect 72882 33567 72894 33570
rect 73490 33567 73502 33570
rect 72882 33521 73502 33567
rect 72882 33518 72894 33521
rect 73490 33518 73502 33521
rect 73554 33518 73566 33570
rect 82126 33506 82178 33518
rect 53454 33458 53506 33470
rect 53454 33394 53506 33406
rect 53790 33458 53842 33470
rect 59726 33458 59778 33470
rect 57362 33406 57374 33458
rect 57426 33406 57438 33458
rect 53790 33394 53842 33406
rect 59726 33394 59778 33406
rect 61406 33458 61458 33470
rect 73502 33458 73554 33470
rect 62066 33406 62078 33458
rect 62130 33406 62142 33458
rect 64194 33406 64206 33458
rect 64258 33406 64270 33458
rect 68562 33406 68574 33458
rect 68626 33406 68638 33458
rect 70466 33406 70478 33458
rect 70530 33406 70542 33458
rect 72594 33406 72606 33458
rect 72658 33406 72670 33458
rect 81106 33406 81118 33458
rect 81170 33406 81182 33458
rect 86482 33406 86494 33458
rect 86546 33406 86558 33458
rect 88610 33406 88622 33458
rect 88674 33406 88686 33458
rect 89506 33406 89518 33458
rect 89570 33406 89582 33458
rect 91634 33406 91646 33458
rect 91698 33406 91710 33458
rect 95330 33406 95342 33458
rect 95394 33406 95406 33458
rect 97458 33406 97470 33458
rect 97522 33406 97534 33458
rect 61406 33394 61458 33406
rect 73502 33394 73554 33406
rect 51662 33346 51714 33358
rect 58382 33346 58434 33358
rect 74286 33346 74338 33358
rect 76302 33346 76354 33358
rect 83918 33346 83970 33358
rect 54450 33294 54462 33346
rect 54514 33294 54526 33346
rect 59154 33294 59166 33346
rect 59218 33294 59230 33346
rect 60386 33294 60398 33346
rect 60450 33294 60462 33346
rect 64978 33294 64990 33346
rect 65042 33294 65054 33346
rect 65762 33294 65774 33346
rect 65826 33294 65838 33346
rect 69682 33294 69694 33346
rect 69746 33294 69758 33346
rect 74722 33294 74734 33346
rect 74786 33294 74798 33346
rect 78306 33294 78318 33346
rect 78370 33294 78382 33346
rect 82786 33294 82798 33346
rect 82850 33294 82862 33346
rect 85810 33294 85822 33346
rect 85874 33294 85886 33346
rect 92418 33294 92430 33346
rect 92482 33294 92494 33346
rect 94546 33294 94558 33346
rect 94610 33294 94622 33346
rect 51662 33282 51714 33294
rect 58382 33282 58434 33294
rect 74286 33282 74338 33294
rect 76302 33282 76354 33294
rect 83918 33282 83970 33294
rect 51326 33234 51378 33246
rect 60622 33234 60674 33246
rect 77310 33234 77362 33246
rect 55234 33182 55246 33234
rect 55298 33182 55310 33234
rect 58930 33182 58942 33234
rect 58994 33182 59006 33234
rect 66434 33182 66446 33234
rect 66498 33182 66510 33234
rect 51326 33170 51378 33182
rect 60622 33170 60674 33182
rect 77310 33170 77362 33182
rect 77646 33234 77698 33246
rect 78978 33182 78990 33234
rect 79042 33182 79054 33234
rect 82898 33182 82910 33234
rect 82962 33182 82974 33234
rect 77646 33170 77698 33182
rect 58046 33122 58098 33134
rect 58046 33058 58098 33070
rect 73054 33122 73106 33134
rect 73054 33058 73106 33070
rect 75742 33122 75794 33134
rect 75742 33058 75794 33070
rect 81790 33122 81842 33134
rect 81790 33058 81842 33070
rect 83582 33122 83634 33134
rect 83582 33058 83634 33070
rect 84366 33122 84418 33134
rect 84366 33058 84418 33070
rect 1344 32954 98560 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 98560 32954
rect 1344 32868 98560 32902
rect 53790 32786 53842 32798
rect 53790 32722 53842 32734
rect 54462 32786 54514 32798
rect 54462 32722 54514 32734
rect 57822 32786 57874 32798
rect 57822 32722 57874 32734
rect 58382 32786 58434 32798
rect 58382 32722 58434 32734
rect 59726 32786 59778 32798
rect 59726 32722 59778 32734
rect 60734 32786 60786 32798
rect 60734 32722 60786 32734
rect 61070 32786 61122 32798
rect 61070 32722 61122 32734
rect 61742 32786 61794 32798
rect 61742 32722 61794 32734
rect 63534 32786 63586 32798
rect 63534 32722 63586 32734
rect 71374 32786 71426 32798
rect 71374 32722 71426 32734
rect 72606 32786 72658 32798
rect 72606 32722 72658 32734
rect 73838 32786 73890 32798
rect 73838 32722 73890 32734
rect 74286 32786 74338 32798
rect 74286 32722 74338 32734
rect 75070 32786 75122 32798
rect 75070 32722 75122 32734
rect 75518 32786 75570 32798
rect 75518 32722 75570 32734
rect 76750 32786 76802 32798
rect 76750 32722 76802 32734
rect 80670 32786 80722 32798
rect 80670 32722 80722 32734
rect 81342 32786 81394 32798
rect 81342 32722 81394 32734
rect 85598 32786 85650 32798
rect 85598 32722 85650 32734
rect 86046 32786 86098 32798
rect 86046 32722 86098 32734
rect 86718 32786 86770 32798
rect 86718 32722 86770 32734
rect 88510 32786 88562 32798
rect 88510 32722 88562 32734
rect 89182 32786 89234 32798
rect 89182 32722 89234 32734
rect 94110 32786 94162 32798
rect 94110 32722 94162 32734
rect 94670 32786 94722 32798
rect 94670 32722 94722 32734
rect 95230 32786 95282 32798
rect 95230 32722 95282 32734
rect 76190 32674 76242 32686
rect 81678 32674 81730 32686
rect 56578 32622 56590 32674
rect 56642 32622 56654 32674
rect 62626 32622 62638 32674
rect 62690 32622 62702 32674
rect 70242 32622 70254 32674
rect 70306 32622 70318 32674
rect 77858 32622 77870 32674
rect 77922 32622 77934 32674
rect 83010 32622 83022 32674
rect 83074 32622 83086 32674
rect 87378 32622 87390 32674
rect 87442 32622 87454 32674
rect 87826 32622 87838 32674
rect 87890 32622 87902 32674
rect 90738 32622 90750 32674
rect 90802 32622 90814 32674
rect 95778 32622 95790 32674
rect 95842 32622 95854 32674
rect 96226 32622 96238 32674
rect 96290 32622 96302 32674
rect 76190 32610 76242 32622
rect 81678 32610 81730 32622
rect 54798 32562 54850 32574
rect 54798 32498 54850 32510
rect 55470 32562 55522 32574
rect 55470 32498 55522 32510
rect 55806 32562 55858 32574
rect 62078 32562 62130 32574
rect 70926 32562 70978 32574
rect 56466 32510 56478 32562
rect 56530 32510 56542 32562
rect 57586 32510 57598 32562
rect 57650 32510 57662 32562
rect 62850 32510 62862 32562
rect 62914 32510 62926 32562
rect 65762 32510 65774 32562
rect 65826 32510 65838 32562
rect 70354 32510 70366 32562
rect 70418 32510 70430 32562
rect 55806 32498 55858 32510
rect 62078 32498 62130 32510
rect 70926 32498 70978 32510
rect 72046 32562 72098 32574
rect 72046 32498 72098 32510
rect 73278 32562 73330 32574
rect 73278 32498 73330 32510
rect 77086 32562 77138 32574
rect 90190 32562 90242 32574
rect 91534 32562 91586 32574
rect 77522 32510 77534 32562
rect 77586 32510 77598 32562
rect 82338 32510 82350 32562
rect 82402 32510 82414 32562
rect 90962 32510 90974 32562
rect 91026 32510 91038 32562
rect 77086 32498 77138 32510
rect 90190 32498 90242 32510
rect 91534 32498 91586 32510
rect 95566 32562 95618 32574
rect 95566 32498 95618 32510
rect 69582 32450 69634 32462
rect 66434 32398 66446 32450
rect 66498 32398 66510 32450
rect 68562 32398 68574 32450
rect 68626 32398 68638 32450
rect 85138 32398 85150 32450
rect 85202 32398 85214 32450
rect 69582 32386 69634 32398
rect 69246 32338 69298 32350
rect 69246 32274 69298 32286
rect 87054 32338 87106 32350
rect 87054 32274 87106 32286
rect 89854 32338 89906 32350
rect 89854 32274 89906 32286
rect 1344 32170 98560 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 98560 32170
rect 1344 32084 98560 32118
rect 57038 31890 57090 31902
rect 57038 31826 57090 31838
rect 57934 31890 57986 31902
rect 57934 31826 57986 31838
rect 61406 31890 61458 31902
rect 61406 31826 61458 31838
rect 68574 31890 68626 31902
rect 68574 31826 68626 31838
rect 70366 31890 70418 31902
rect 76414 31890 76466 31902
rect 71586 31838 71598 31890
rect 71650 31838 71662 31890
rect 73714 31838 73726 31890
rect 73778 31838 73790 31890
rect 70366 31826 70418 31838
rect 76414 31826 76466 31838
rect 86942 31890 86994 31902
rect 86942 31826 86994 31838
rect 89294 31890 89346 31902
rect 89294 31826 89346 31838
rect 55918 31778 55970 31790
rect 55918 31714 55970 31726
rect 67006 31778 67058 31790
rect 67006 31714 67058 31726
rect 68014 31778 68066 31790
rect 70802 31726 70814 31778
rect 70866 31726 70878 31778
rect 89842 31726 89854 31778
rect 89906 31726 89918 31778
rect 68014 31714 68066 31726
rect 55582 31666 55634 31678
rect 55582 31602 55634 31614
rect 66670 31666 66722 31678
rect 66670 31602 66722 31614
rect 67678 31666 67730 31678
rect 67678 31602 67730 31614
rect 69358 31666 69410 31678
rect 69358 31602 69410 31614
rect 69694 31666 69746 31678
rect 69694 31602 69746 31614
rect 84142 31666 84194 31678
rect 84142 31602 84194 31614
rect 90078 31666 90130 31678
rect 90078 31602 90130 31614
rect 57374 31554 57426 31566
rect 57374 31490 57426 31502
rect 83806 31554 83858 31566
rect 83806 31490 83858 31502
rect 1344 31386 98560 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 98560 31386
rect 1344 31300 98560 31334
rect 70590 31218 70642 31230
rect 70590 31154 70642 31166
rect 83906 31054 83918 31106
rect 83970 31054 83982 31106
rect 83122 30942 83134 30994
rect 83186 30942 83198 30994
rect 69022 30882 69074 30894
rect 86034 30830 86046 30882
rect 86098 30830 86110 30882
rect 69022 30818 69074 30830
rect 1344 30602 98560 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 98560 30602
rect 1344 30516 98560 30550
rect 1344 29818 98560 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 98560 29818
rect 1344 29732 98560 29766
rect 83694 29650 83746 29662
rect 83694 29586 83746 29598
rect 84254 29650 84306 29662
rect 84254 29586 84306 29598
rect 85138 29486 85150 29538
rect 85202 29486 85214 29538
rect 83246 29426 83298 29438
rect 83246 29362 83298 29374
rect 84590 29426 84642 29438
rect 85362 29374 85374 29426
rect 85426 29374 85438 29426
rect 84590 29362 84642 29374
rect 1344 29034 98560 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 98560 29034
rect 1344 28948 98560 28982
rect 1344 28250 98560 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 98560 28250
rect 1344 28164 98560 28198
rect 1344 27466 98560 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 98560 27466
rect 1344 27380 98560 27414
rect 1344 26682 98560 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 98560 26682
rect 1344 26596 98560 26630
rect 1344 25898 98560 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 98560 25898
rect 1344 25812 98560 25846
rect 95230 25394 95282 25406
rect 95230 25330 95282 25342
rect 94894 25282 94946 25294
rect 94894 25218 94946 25230
rect 95790 25282 95842 25294
rect 95790 25218 95842 25230
rect 1344 25114 98560 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 98560 25114
rect 1344 25028 98560 25062
rect 1344 24330 98560 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 98560 24330
rect 1344 24244 98560 24278
rect 1344 23546 98560 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 98560 23546
rect 1344 23460 98560 23494
rect 1344 22762 98560 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 98560 22762
rect 1344 22676 98560 22710
rect 1344 21978 98560 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 98560 21978
rect 1344 21892 98560 21926
rect 1344 21194 98560 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 98560 21194
rect 1344 21108 98560 21142
rect 1344 20410 98560 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 98560 20410
rect 1344 20324 98560 20358
rect 1344 19626 98560 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 98560 19626
rect 1344 19540 98560 19574
rect 1344 18842 98560 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 98560 18842
rect 1344 18756 98560 18790
rect 1344 18058 98560 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 98560 18058
rect 1344 17972 98560 18006
rect 1344 17274 98560 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 98560 17274
rect 1344 17188 98560 17222
rect 1344 16490 98560 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 98560 16490
rect 1344 16404 98560 16438
rect 1344 15706 98560 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 98560 15706
rect 1344 15620 98560 15654
rect 1344 14922 98560 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 98560 14922
rect 1344 14836 98560 14870
rect 1344 14138 98560 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 98560 14138
rect 1344 14052 98560 14086
rect 1344 13354 98560 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 98560 13354
rect 1344 13268 98560 13302
rect 1822 12850 1874 12862
rect 1822 12786 1874 12798
rect 2158 12738 2210 12750
rect 2158 12674 2210 12686
rect 1344 12570 98560 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 98560 12570
rect 1344 12484 98560 12518
rect 1822 12402 1874 12414
rect 1822 12338 1874 12350
rect 1344 11786 98560 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 98560 11786
rect 1344 11700 98560 11734
rect 1344 11002 98560 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 98560 11002
rect 1344 10916 98560 10950
rect 1344 10218 98560 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 98560 10218
rect 1344 10132 98560 10166
rect 1344 9434 98560 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 98560 9434
rect 1344 9348 98560 9382
rect 1344 8650 98560 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 98560 8650
rect 1344 8564 98560 8598
rect 1344 7866 98560 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 98560 7866
rect 1344 7780 98560 7814
rect 1344 7082 98560 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 98560 7082
rect 1344 6996 98560 7030
rect 1344 6298 98560 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 98560 6298
rect 1344 6212 98560 6246
rect 1344 5514 98560 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 98560 5514
rect 1344 5428 98560 5462
rect 1344 4730 98560 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 98560 4730
rect 1344 4644 98560 4678
rect 1344 3946 98560 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 98560 3946
rect 1344 3860 98560 3894
rect 6190 3442 6242 3454
rect 6190 3378 6242 3390
rect 6638 3442 6690 3454
rect 6638 3378 6690 3390
rect 18622 3442 18674 3454
rect 18622 3378 18674 3390
rect 19070 3442 19122 3454
rect 19070 3378 19122 3390
rect 31054 3442 31106 3454
rect 31054 3378 31106 3390
rect 31502 3442 31554 3454
rect 31502 3378 31554 3390
rect 44270 3442 44322 3454
rect 44270 3378 44322 3390
rect 44942 3442 44994 3454
rect 44942 3378 44994 3390
rect 56030 3442 56082 3454
rect 56030 3378 56082 3390
rect 56702 3442 56754 3454
rect 56702 3378 56754 3390
rect 67790 3442 67842 3454
rect 67790 3378 67842 3390
rect 68798 3442 68850 3454
rect 68798 3378 68850 3390
rect 80782 3442 80834 3454
rect 80782 3378 80834 3390
rect 81230 3442 81282 3454
rect 81230 3378 81282 3390
rect 93214 3442 93266 3454
rect 93214 3378 93266 3390
rect 93998 3442 94050 3454
rect 93998 3378 94050 3390
rect 6974 3330 7026 3342
rect 6974 3266 7026 3278
rect 19406 3330 19458 3342
rect 19406 3266 19458 3278
rect 31838 3330 31890 3342
rect 31838 3266 31890 3278
rect 45278 3330 45330 3342
rect 45278 3266 45330 3278
rect 57038 3330 57090 3342
rect 57038 3266 57090 3278
rect 69134 3330 69186 3342
rect 69134 3266 69186 3278
rect 81566 3330 81618 3342
rect 81566 3266 81618 3278
rect 93662 3330 93714 3342
rect 93662 3266 93714 3278
rect 1344 3162 98560 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 98560 3162
rect 1344 3076 98560 3110
<< via1 >>
rect 43710 96574 43762 96626
rect 45054 96574 45106 96626
rect 56142 96574 56194 96626
rect 56814 96574 56866 96626
rect 4478 96406 4530 96458
rect 4582 96406 4634 96458
rect 4686 96406 4738 96458
rect 35198 96406 35250 96458
rect 35302 96406 35354 96458
rect 35406 96406 35458 96458
rect 65918 96406 65970 96458
rect 66022 96406 66074 96458
rect 66126 96406 66178 96458
rect 96638 96406 96690 96458
rect 96742 96406 96794 96458
rect 96846 96406 96898 96458
rect 6750 96126 6802 96178
rect 19182 96126 19234 96178
rect 31278 96126 31330 96178
rect 45054 96126 45106 96178
rect 56814 96126 56866 96178
rect 68910 96126 68962 96178
rect 81342 96126 81394 96178
rect 94334 96126 94386 96178
rect 7870 96014 7922 96066
rect 8318 96014 8370 96066
rect 20302 96014 20354 96066
rect 32174 96014 32226 96066
rect 45950 96014 46002 96066
rect 57710 96014 57762 96066
rect 58382 96014 58434 96066
rect 70030 96014 70082 96066
rect 82350 96014 82402 96066
rect 93102 96014 93154 96066
rect 93886 96014 93938 96066
rect 21310 95790 21362 95842
rect 33070 95790 33122 95842
rect 46622 95790 46674 95842
rect 70478 95790 70530 95842
rect 82910 95790 82962 95842
rect 19838 95622 19890 95674
rect 19942 95622 19994 95674
rect 20046 95622 20098 95674
rect 50558 95622 50610 95674
rect 50662 95622 50714 95674
rect 50766 95622 50818 95674
rect 81278 95622 81330 95674
rect 81382 95622 81434 95674
rect 81486 95622 81538 95674
rect 4478 94838 4530 94890
rect 4582 94838 4634 94890
rect 4686 94838 4738 94890
rect 35198 94838 35250 94890
rect 35302 94838 35354 94890
rect 35406 94838 35458 94890
rect 65918 94838 65970 94890
rect 66022 94838 66074 94890
rect 66126 94838 66178 94890
rect 96638 94838 96690 94890
rect 96742 94838 96794 94890
rect 96846 94838 96898 94890
rect 19838 94054 19890 94106
rect 19942 94054 19994 94106
rect 20046 94054 20098 94106
rect 50558 94054 50610 94106
rect 50662 94054 50714 94106
rect 50766 94054 50818 94106
rect 81278 94054 81330 94106
rect 81382 94054 81434 94106
rect 81486 94054 81538 94106
rect 4478 93270 4530 93322
rect 4582 93270 4634 93322
rect 4686 93270 4738 93322
rect 35198 93270 35250 93322
rect 35302 93270 35354 93322
rect 35406 93270 35458 93322
rect 65918 93270 65970 93322
rect 66022 93270 66074 93322
rect 66126 93270 66178 93322
rect 96638 93270 96690 93322
rect 96742 93270 96794 93322
rect 96846 93270 96898 93322
rect 19838 92486 19890 92538
rect 19942 92486 19994 92538
rect 20046 92486 20098 92538
rect 50558 92486 50610 92538
rect 50662 92486 50714 92538
rect 50766 92486 50818 92538
rect 81278 92486 81330 92538
rect 81382 92486 81434 92538
rect 81486 92486 81538 92538
rect 4478 91702 4530 91754
rect 4582 91702 4634 91754
rect 4686 91702 4738 91754
rect 35198 91702 35250 91754
rect 35302 91702 35354 91754
rect 35406 91702 35458 91754
rect 65918 91702 65970 91754
rect 66022 91702 66074 91754
rect 66126 91702 66178 91754
rect 96638 91702 96690 91754
rect 96742 91702 96794 91754
rect 96846 91702 96898 91754
rect 19838 90918 19890 90970
rect 19942 90918 19994 90970
rect 20046 90918 20098 90970
rect 50558 90918 50610 90970
rect 50662 90918 50714 90970
rect 50766 90918 50818 90970
rect 81278 90918 81330 90970
rect 81382 90918 81434 90970
rect 81486 90918 81538 90970
rect 4478 90134 4530 90186
rect 4582 90134 4634 90186
rect 4686 90134 4738 90186
rect 35198 90134 35250 90186
rect 35302 90134 35354 90186
rect 35406 90134 35458 90186
rect 65918 90134 65970 90186
rect 66022 90134 66074 90186
rect 66126 90134 66178 90186
rect 96638 90134 96690 90186
rect 96742 90134 96794 90186
rect 96846 90134 96898 90186
rect 19838 89350 19890 89402
rect 19942 89350 19994 89402
rect 20046 89350 20098 89402
rect 50558 89350 50610 89402
rect 50662 89350 50714 89402
rect 50766 89350 50818 89402
rect 81278 89350 81330 89402
rect 81382 89350 81434 89402
rect 81486 89350 81538 89402
rect 68238 88958 68290 89010
rect 90862 88958 90914 89010
rect 63086 88846 63138 88898
rect 63534 88846 63586 88898
rect 68910 88846 68962 88898
rect 71038 88846 71090 88898
rect 71598 88846 71650 88898
rect 91646 88846 91698 88898
rect 93774 88846 93826 88898
rect 4478 88566 4530 88618
rect 4582 88566 4634 88618
rect 4686 88566 4738 88618
rect 35198 88566 35250 88618
rect 35302 88566 35354 88618
rect 35406 88566 35458 88618
rect 65918 88566 65970 88618
rect 66022 88566 66074 88618
rect 66126 88566 66178 88618
rect 96638 88566 96690 88618
rect 96742 88566 96794 88618
rect 96846 88566 96898 88618
rect 3278 88286 3330 88338
rect 61854 88174 61906 88226
rect 62526 88174 62578 88226
rect 1934 88062 1986 88114
rect 57710 88062 57762 88114
rect 62638 88062 62690 88114
rect 63534 88062 63586 88114
rect 54798 87950 54850 88002
rect 57374 87950 57426 88002
rect 59614 87950 59666 88002
rect 60622 87950 60674 88002
rect 61518 87950 61570 88002
rect 63870 87950 63922 88002
rect 64430 87950 64482 88002
rect 70478 87950 70530 88002
rect 71038 87950 71090 88002
rect 19838 87782 19890 87834
rect 19942 87782 19994 87834
rect 20046 87782 20098 87834
rect 50558 87782 50610 87834
rect 50662 87782 50714 87834
rect 50766 87782 50818 87834
rect 81278 87782 81330 87834
rect 81382 87782 81434 87834
rect 81486 87782 81538 87834
rect 58046 87614 58098 87666
rect 54350 87502 54402 87554
rect 59166 87502 59218 87554
rect 64318 87502 64370 87554
rect 72270 87502 72322 87554
rect 87278 87502 87330 87554
rect 89518 87502 89570 87554
rect 1710 87390 1762 87442
rect 54238 87390 54290 87442
rect 55582 87390 55634 87442
rect 56030 87390 56082 87442
rect 59054 87390 59106 87442
rect 59950 87390 60002 87442
rect 64542 87390 64594 87442
rect 65326 87390 65378 87442
rect 67454 87390 67506 87442
rect 70702 87390 70754 87442
rect 72494 87390 72546 87442
rect 87054 87390 87106 87442
rect 94558 87390 94610 87442
rect 95118 87390 95170 87442
rect 55022 87278 55074 87330
rect 57486 87278 57538 87330
rect 60622 87278 60674 87330
rect 62750 87278 62802 87330
rect 68126 87278 68178 87330
rect 70254 87278 70306 87330
rect 73278 87278 73330 87330
rect 73726 87278 73778 87330
rect 74510 87278 74562 87330
rect 75070 87278 75122 87330
rect 75518 87278 75570 87330
rect 53230 87166 53282 87218
rect 53566 87166 53618 87218
rect 58382 87166 58434 87218
rect 63422 87166 63474 87218
rect 63758 87166 63810 87218
rect 71374 87166 71426 87218
rect 71710 87166 71762 87218
rect 4478 86998 4530 87050
rect 4582 86998 4634 87050
rect 4686 86998 4738 87050
rect 35198 86998 35250 87050
rect 35302 86998 35354 87050
rect 35406 86998 35458 87050
rect 65918 86998 65970 87050
rect 66022 86998 66074 87050
rect 66126 86998 66178 87050
rect 96638 86998 96690 87050
rect 96742 86998 96794 87050
rect 96846 86998 96898 87050
rect 81790 86830 81842 86882
rect 87614 86830 87666 86882
rect 57150 86718 57202 86770
rect 59278 86718 59330 86770
rect 60622 86718 60674 86770
rect 62190 86718 62242 86770
rect 65774 86718 65826 86770
rect 73166 86718 73218 86770
rect 74734 86718 74786 86770
rect 52558 86606 52610 86658
rect 53902 86606 53954 86658
rect 54686 86606 54738 86658
rect 55582 86606 55634 86658
rect 56478 86606 56530 86658
rect 60062 86606 60114 86658
rect 61630 86606 61682 86658
rect 62974 86606 63026 86658
rect 69806 86606 69858 86658
rect 71710 86606 71762 86658
rect 73726 86606 73778 86658
rect 74398 86606 74450 86658
rect 77870 86606 77922 86658
rect 87950 86606 88002 86658
rect 54462 86494 54514 86546
rect 61406 86494 61458 86546
rect 63646 86494 63698 86546
rect 68238 86494 68290 86546
rect 68574 86494 68626 86546
rect 70142 86494 70194 86546
rect 70366 86494 70418 86546
rect 71374 86494 71426 86546
rect 71934 86494 71986 86546
rect 72270 86494 72322 86546
rect 75742 86494 75794 86546
rect 81902 86494 81954 86546
rect 82462 86494 82514 86546
rect 86494 86494 86546 86546
rect 88174 86494 88226 86546
rect 88734 86494 88786 86546
rect 91534 86494 91586 86546
rect 91870 86494 91922 86546
rect 95566 86494 95618 86546
rect 52222 86382 52274 86434
rect 53566 86382 53618 86434
rect 55358 86382 55410 86434
rect 59838 86382 59890 86434
rect 66334 86382 66386 86434
rect 66670 86382 66722 86434
rect 69470 86382 69522 86434
rect 75406 86382 75458 86434
rect 76526 86382 76578 86434
rect 77310 86382 77362 86434
rect 78094 86382 78146 86434
rect 78654 86382 78706 86434
rect 79662 86382 79714 86434
rect 81230 86382 81282 86434
rect 81790 86382 81842 86434
rect 82574 86382 82626 86434
rect 82798 86382 82850 86434
rect 83134 86382 83186 86434
rect 86158 86382 86210 86434
rect 87054 86382 87106 86434
rect 89294 86382 89346 86434
rect 95902 86382 95954 86434
rect 19838 86214 19890 86266
rect 19942 86214 19994 86266
rect 20046 86214 20098 86266
rect 50558 86214 50610 86266
rect 50662 86214 50714 86266
rect 50766 86214 50818 86266
rect 81278 86214 81330 86266
rect 81382 86214 81434 86266
rect 81486 86214 81538 86266
rect 55470 86046 55522 86098
rect 72718 86046 72770 86098
rect 73390 86046 73442 86098
rect 79214 86046 79266 86098
rect 56590 85934 56642 85986
rect 58270 85934 58322 85986
rect 75294 85934 75346 85986
rect 78206 85934 78258 85986
rect 78654 85934 78706 85986
rect 87726 85934 87778 85986
rect 95902 85934 95954 85986
rect 51214 85822 51266 85874
rect 56478 85822 56530 85874
rect 57598 85822 57650 85874
rect 63086 85822 63138 85874
rect 63870 85822 63922 85874
rect 66446 85822 66498 85874
rect 74622 85822 74674 85874
rect 84254 85822 84306 85874
rect 88398 85822 88450 85874
rect 93550 85822 93602 85874
rect 95566 85822 95618 85874
rect 51886 85710 51938 85762
rect 54014 85710 54066 85762
rect 54574 85710 54626 85762
rect 55806 85710 55858 85762
rect 60398 85710 60450 85762
rect 60958 85710 61010 85762
rect 64318 85710 64370 85762
rect 65438 85710 65490 85762
rect 69470 85710 69522 85762
rect 71710 85710 71762 85762
rect 73838 85710 73890 85762
rect 77422 85710 77474 85762
rect 78878 85710 78930 85762
rect 79774 85710 79826 85762
rect 80446 85710 80498 85762
rect 81342 85710 81394 85762
rect 83470 85710 83522 85762
rect 84814 85710 84866 85762
rect 85598 85710 85650 85762
rect 89182 85710 89234 85762
rect 90638 85710 90690 85762
rect 92766 85710 92818 85762
rect 4478 85430 4530 85482
rect 4582 85430 4634 85482
rect 4686 85430 4738 85482
rect 35198 85430 35250 85482
rect 35302 85430 35354 85482
rect 35406 85430 35458 85482
rect 65918 85430 65970 85482
rect 66022 85430 66074 85482
rect 66126 85430 66178 85482
rect 96638 85430 96690 85482
rect 96742 85430 96794 85482
rect 96846 85430 96898 85482
rect 59390 85262 59442 85314
rect 59726 85262 59778 85314
rect 74958 85262 75010 85314
rect 75294 85262 75346 85314
rect 88846 85262 88898 85314
rect 91198 85262 91250 85314
rect 55134 85150 55186 85202
rect 57262 85150 57314 85202
rect 57710 85150 57762 85202
rect 60286 85150 60338 85202
rect 62638 85150 62690 85202
rect 64766 85150 64818 85202
rect 72270 85150 72322 85202
rect 73166 85150 73218 85202
rect 86046 85150 86098 85202
rect 88174 85150 88226 85202
rect 89182 85150 89234 85202
rect 95678 85150 95730 85202
rect 97806 85150 97858 85202
rect 52558 85038 52610 85090
rect 54462 85038 54514 85090
rect 61518 85038 61570 85090
rect 65550 85038 65602 85090
rect 66558 85038 66610 85090
rect 67118 85038 67170 85090
rect 68350 85038 68402 85090
rect 69470 85038 69522 85090
rect 74062 85038 74114 85090
rect 82574 85038 82626 85090
rect 85374 85038 85426 85090
rect 89630 85038 89682 85090
rect 91534 85038 91586 85090
rect 92206 85038 92258 85090
rect 93438 85038 93490 85090
rect 94894 85038 94946 85090
rect 52222 84926 52274 84978
rect 58718 84926 58770 84978
rect 59054 84926 59106 84978
rect 61742 84926 61794 84978
rect 67230 84926 67282 84978
rect 70142 84926 70194 84978
rect 75630 84926 75682 84978
rect 76078 84926 76130 84978
rect 78766 84926 78818 84978
rect 89742 84926 89794 84978
rect 92318 84926 92370 84978
rect 93214 84926 93266 84978
rect 53790 84814 53842 84866
rect 66222 84814 66274 84866
rect 68014 84814 68066 84866
rect 72830 84814 72882 84866
rect 74286 84814 74338 84866
rect 83022 84814 83074 84866
rect 83470 84814 83522 84866
rect 90526 84814 90578 84866
rect 94446 84814 94498 84866
rect 19838 84646 19890 84698
rect 19942 84646 19994 84698
rect 20046 84646 20098 84698
rect 50558 84646 50610 84698
rect 50662 84646 50714 84698
rect 50766 84646 50818 84698
rect 81278 84646 81330 84698
rect 81382 84646 81434 84698
rect 81486 84646 81538 84698
rect 65774 84478 65826 84530
rect 90526 84478 90578 84530
rect 95230 84478 95282 84530
rect 51774 84366 51826 84418
rect 60622 84366 60674 84418
rect 67118 84366 67170 84418
rect 71038 84366 71090 84418
rect 74286 84366 74338 84418
rect 78094 84366 78146 84418
rect 84926 84366 84978 84418
rect 87726 84366 87778 84418
rect 89294 84366 89346 84418
rect 95790 84366 95842 84418
rect 96350 84366 96402 84418
rect 51102 84254 51154 84306
rect 58830 84254 58882 84306
rect 64318 84254 64370 84306
rect 66334 84254 66386 84306
rect 71262 84254 71314 84306
rect 71934 84254 71986 84306
rect 72494 84254 72546 84306
rect 73614 84254 73666 84306
rect 77422 84254 77474 84306
rect 81454 84254 81506 84306
rect 85038 84254 85090 84306
rect 88510 84254 88562 84306
rect 89518 84254 89570 84306
rect 90190 84254 90242 84306
rect 94446 84254 94498 84306
rect 95566 84254 95618 84306
rect 53902 84142 53954 84194
rect 54462 84142 54514 84194
rect 54798 84142 54850 84194
rect 57374 84142 57426 84194
rect 69246 84142 69298 84194
rect 76414 84142 76466 84194
rect 80222 84142 80274 84194
rect 82126 84142 82178 84194
rect 84254 84142 84306 84194
rect 85598 84142 85650 84194
rect 90974 84142 91026 84194
rect 91534 84142 91586 84194
rect 93662 84142 93714 84194
rect 70142 84030 70194 84082
rect 70478 84030 70530 84082
rect 84926 84030 84978 84082
rect 4478 83862 4530 83914
rect 4582 83862 4634 83914
rect 4686 83862 4738 83914
rect 35198 83862 35250 83914
rect 35302 83862 35354 83914
rect 35406 83862 35458 83914
rect 65918 83862 65970 83914
rect 66022 83862 66074 83914
rect 66126 83862 66178 83914
rect 96638 83862 96690 83914
rect 96742 83862 96794 83914
rect 96846 83862 96898 83914
rect 63422 83694 63474 83746
rect 74286 83694 74338 83746
rect 74622 83694 74674 83746
rect 83694 83694 83746 83746
rect 88286 83694 88338 83746
rect 88622 83694 88674 83746
rect 91198 83694 91250 83746
rect 65102 83582 65154 83634
rect 67678 83582 67730 83634
rect 79550 83582 79602 83634
rect 83022 83582 83074 83634
rect 90526 83582 90578 83634
rect 94334 83582 94386 83634
rect 95678 83582 95730 83634
rect 97806 83582 97858 83634
rect 53678 83470 53730 83522
rect 57934 83470 57986 83522
rect 63758 83470 63810 83522
rect 64430 83470 64482 83522
rect 69694 83470 69746 83522
rect 70590 83470 70642 83522
rect 72718 83470 72770 83522
rect 73166 83470 73218 83522
rect 77534 83470 77586 83522
rect 78206 83470 78258 83522
rect 80222 83470 80274 83522
rect 91534 83470 91586 83522
rect 92206 83470 92258 83522
rect 93326 83470 93378 83522
rect 94894 83470 94946 83522
rect 54462 83358 54514 83410
rect 64542 83358 64594 83410
rect 69358 83358 69410 83410
rect 70254 83358 70306 83410
rect 74958 83358 75010 83410
rect 75406 83358 75458 83410
rect 76414 83358 76466 83410
rect 77422 83358 77474 83410
rect 78542 83358 78594 83410
rect 80894 83358 80946 83410
rect 83582 83358 83634 83410
rect 88846 83358 88898 83410
rect 89406 83358 89458 83410
rect 92318 83358 92370 83410
rect 93550 83358 93602 83410
rect 52670 83246 52722 83298
rect 53342 83246 53394 83298
rect 53566 83246 53618 83298
rect 54126 83246 54178 83298
rect 54350 83246 54402 83298
rect 54910 83246 54962 83298
rect 56926 83246 56978 83298
rect 58158 83246 58210 83298
rect 71598 83246 71650 83298
rect 73614 83246 73666 83298
rect 76078 83246 76130 83298
rect 79214 83246 79266 83298
rect 83694 83246 83746 83298
rect 84366 83246 84418 83298
rect 85262 83246 85314 83298
rect 85710 83246 85762 83298
rect 87614 83246 87666 83298
rect 19838 83078 19890 83130
rect 19942 83078 19994 83130
rect 20046 83078 20098 83130
rect 50558 83078 50610 83130
rect 50662 83078 50714 83130
rect 50766 83078 50818 83130
rect 81278 83078 81330 83130
rect 81382 83078 81434 83130
rect 81486 83078 81538 83130
rect 60846 82910 60898 82962
rect 63422 82910 63474 82962
rect 74846 82910 74898 82962
rect 78766 82910 78818 82962
rect 80446 82910 80498 82962
rect 58270 82798 58322 82850
rect 61630 82798 61682 82850
rect 63758 82798 63810 82850
rect 76190 82798 76242 82850
rect 82686 82798 82738 82850
rect 52894 82686 52946 82738
rect 57598 82686 57650 82738
rect 61966 82686 62018 82738
rect 75518 82686 75570 82738
rect 80334 82686 80386 82738
rect 82014 82686 82066 82738
rect 92654 82686 92706 82738
rect 54126 82574 54178 82626
rect 60398 82574 60450 82626
rect 69470 82574 69522 82626
rect 69918 82574 69970 82626
rect 73838 82574 73890 82626
rect 78318 82574 78370 82626
rect 81454 82574 81506 82626
rect 84814 82574 84866 82626
rect 85262 82574 85314 82626
rect 85822 82574 85874 82626
rect 86158 82574 86210 82626
rect 86606 82574 86658 82626
rect 90638 82574 90690 82626
rect 94894 82574 94946 82626
rect 80446 82462 80498 82514
rect 85710 82462 85762 82514
rect 86718 82462 86770 82514
rect 4478 82294 4530 82346
rect 4582 82294 4634 82346
rect 4686 82294 4738 82346
rect 35198 82294 35250 82346
rect 35302 82294 35354 82346
rect 35406 82294 35458 82346
rect 65918 82294 65970 82346
rect 66022 82294 66074 82346
rect 66126 82294 66178 82346
rect 96638 82294 96690 82346
rect 96742 82294 96794 82346
rect 96846 82294 96898 82346
rect 58606 82126 58658 82178
rect 62302 82126 62354 82178
rect 93326 82126 93378 82178
rect 95230 82126 95282 82178
rect 52670 82014 52722 82066
rect 57038 82014 57090 82066
rect 63982 82014 64034 82066
rect 73278 82014 73330 82066
rect 75406 82014 75458 82066
rect 77870 82014 77922 82066
rect 97358 82014 97410 82066
rect 49758 81902 49810 81954
rect 54126 81902 54178 81954
rect 58942 81902 58994 81954
rect 59726 81902 59778 81954
rect 62638 81902 62690 81954
rect 63422 81902 63474 81954
rect 81118 81902 81170 81954
rect 81454 81902 81506 81954
rect 82686 81902 82738 81954
rect 83022 81902 83074 81954
rect 83918 81902 83970 81954
rect 86718 81902 86770 81954
rect 93662 81902 93714 81954
rect 95566 81902 95618 81954
rect 96238 81902 96290 81954
rect 50542 81790 50594 81842
rect 54910 81790 54962 81842
rect 59502 81790 59554 81842
rect 63198 81790 63250 81842
rect 68014 81790 68066 81842
rect 72830 81790 72882 81842
rect 83582 81790 83634 81842
rect 87614 81790 87666 81842
rect 93886 81790 93938 81842
rect 94222 81790 94274 81842
rect 96350 81790 96402 81842
rect 53342 81678 53394 81730
rect 60286 81678 60338 81730
rect 64430 81678 64482 81730
rect 68126 81678 68178 81730
rect 68350 81678 68402 81730
rect 69806 81678 69858 81730
rect 70366 81678 70418 81730
rect 73838 81678 73890 81730
rect 74286 81678 74338 81730
rect 74846 81678 74898 81730
rect 76526 81678 76578 81730
rect 77310 81678 77362 81730
rect 80670 81678 80722 81730
rect 81342 81678 81394 81730
rect 82014 81678 82066 81730
rect 82910 81678 82962 81730
rect 83694 81678 83746 81730
rect 84366 81678 84418 81730
rect 90974 81678 91026 81730
rect 92430 81678 92482 81730
rect 96910 81678 96962 81730
rect 97806 81678 97858 81730
rect 19838 81510 19890 81562
rect 19942 81510 19994 81562
rect 20046 81510 20098 81562
rect 50558 81510 50610 81562
rect 50662 81510 50714 81562
rect 50766 81510 50818 81562
rect 81278 81510 81330 81562
rect 81382 81510 81434 81562
rect 81486 81510 81538 81562
rect 50766 81342 50818 81394
rect 56590 81342 56642 81394
rect 69694 81342 69746 81394
rect 73838 81342 73890 81394
rect 74510 81342 74562 81394
rect 75070 81342 75122 81394
rect 80558 81342 80610 81394
rect 92206 81342 92258 81394
rect 50206 81230 50258 81282
rect 50318 81230 50370 81282
rect 50990 81230 51042 81282
rect 52446 81230 52498 81282
rect 55246 81230 55298 81282
rect 56030 81230 56082 81282
rect 61294 81230 61346 81282
rect 63982 81230 64034 81282
rect 68462 81230 68514 81282
rect 81454 81230 81506 81282
rect 82350 81230 82402 81282
rect 83134 81230 83186 81282
rect 83246 81230 83298 81282
rect 85262 81230 85314 81282
rect 86270 81230 86322 81282
rect 93550 81230 93602 81282
rect 93774 81230 93826 81282
rect 95790 81230 95842 81282
rect 96126 81230 96178 81282
rect 51102 81118 51154 81170
rect 51662 81118 51714 81170
rect 55022 81118 55074 81170
rect 55358 81118 55410 81170
rect 55806 81118 55858 81170
rect 56142 81118 56194 81170
rect 60622 81118 60674 81170
rect 64206 81118 64258 81170
rect 69246 81118 69298 81170
rect 71486 81118 71538 81170
rect 72606 81118 72658 81170
rect 73502 81118 73554 81170
rect 74286 81118 74338 81170
rect 74622 81118 74674 81170
rect 80110 81118 80162 81170
rect 81566 81118 81618 81170
rect 82126 81118 82178 81170
rect 82462 81118 82514 81170
rect 82910 81118 82962 81170
rect 85710 81118 85762 81170
rect 86046 81118 86098 81170
rect 86830 81118 86882 81170
rect 87502 81118 87554 81170
rect 88398 81118 88450 81170
rect 54574 81006 54626 81058
rect 57374 81006 57426 81058
rect 63422 81006 63474 81058
rect 66334 81006 66386 81058
rect 70142 81006 70194 81058
rect 70590 81006 70642 81058
rect 71150 81006 71202 81058
rect 72046 81006 72098 81058
rect 83694 81006 83746 81058
rect 84142 81006 84194 81058
rect 84590 81006 84642 81058
rect 93214 81006 93266 81058
rect 94670 81006 94722 81058
rect 95566 81006 95618 81058
rect 97246 81006 97298 81058
rect 50206 80894 50258 80946
rect 71150 80894 71202 80946
rect 71598 80894 71650 80946
rect 72046 80894 72098 80946
rect 81454 80894 81506 80946
rect 92878 80894 92930 80946
rect 95230 80894 95282 80946
rect 4478 80726 4530 80778
rect 4582 80726 4634 80778
rect 4686 80726 4738 80778
rect 35198 80726 35250 80778
rect 35302 80726 35354 80778
rect 35406 80726 35458 80778
rect 65918 80726 65970 80778
rect 66022 80726 66074 80778
rect 66126 80726 66178 80778
rect 96638 80726 96690 80778
rect 96742 80726 96794 80778
rect 96846 80726 96898 80778
rect 83582 80558 83634 80610
rect 85710 80558 85762 80610
rect 86494 80558 86546 80610
rect 52334 80446 52386 80498
rect 54238 80446 54290 80498
rect 56366 80446 56418 80498
rect 61406 80446 61458 80498
rect 63534 80446 63586 80498
rect 68574 80446 68626 80498
rect 74510 80446 74562 80498
rect 79550 80446 79602 80498
rect 81678 80446 81730 80498
rect 85598 80446 85650 80498
rect 86046 80446 86098 80498
rect 86494 80446 86546 80498
rect 88510 80446 88562 80498
rect 93102 80446 93154 80498
rect 93550 80446 93602 80498
rect 97806 80446 97858 80498
rect 49534 80334 49586 80386
rect 53454 80334 53506 80386
rect 56814 80334 56866 80386
rect 57150 80334 57202 80386
rect 57598 80334 57650 80386
rect 64318 80334 64370 80386
rect 65774 80334 65826 80386
rect 70030 80334 70082 80386
rect 70366 80334 70418 80386
rect 71710 80334 71762 80386
rect 75294 80334 75346 80386
rect 78878 80334 78930 80386
rect 82910 80334 82962 80386
rect 84254 80334 84306 80386
rect 92430 80334 92482 80386
rect 94894 80334 94946 80386
rect 50206 80222 50258 80274
rect 57038 80222 57090 80274
rect 66446 80222 66498 80274
rect 69470 80222 69522 80274
rect 69582 80222 69634 80274
rect 70814 80222 70866 80274
rect 72382 80222 72434 80274
rect 74958 80222 75010 80274
rect 75182 80222 75234 80274
rect 83582 80222 83634 80274
rect 83694 80222 83746 80274
rect 94334 80222 94386 80274
rect 95678 80222 95730 80274
rect 64766 80110 64818 80162
rect 69246 80110 69298 80162
rect 70254 80110 70306 80162
rect 75742 80110 75794 80162
rect 76190 80110 76242 80162
rect 82238 80110 82290 80162
rect 82574 80110 82626 80162
rect 82798 80110 82850 80162
rect 84366 80110 84418 80162
rect 84590 80110 84642 80162
rect 85150 80110 85202 80162
rect 19838 79942 19890 79994
rect 19942 79942 19994 79994
rect 20046 79942 20098 79994
rect 50558 79942 50610 79994
rect 50662 79942 50714 79994
rect 50766 79942 50818 79994
rect 81278 79942 81330 79994
rect 81382 79942 81434 79994
rect 81486 79942 81538 79994
rect 52894 79774 52946 79826
rect 53118 79774 53170 79826
rect 53678 79774 53730 79826
rect 54350 79774 54402 79826
rect 55134 79774 55186 79826
rect 55918 79774 55970 79826
rect 56702 79774 56754 79826
rect 63646 79774 63698 79826
rect 64318 79774 64370 79826
rect 70814 79774 70866 79826
rect 71374 79774 71426 79826
rect 72270 79774 72322 79826
rect 80446 79774 80498 79826
rect 84702 79774 84754 79826
rect 89182 79774 89234 79826
rect 89630 79774 89682 79826
rect 97246 79774 97298 79826
rect 50318 79662 50370 79714
rect 53230 79662 53282 79714
rect 54574 79662 54626 79714
rect 55358 79662 55410 79714
rect 55470 79662 55522 79714
rect 57486 79662 57538 79714
rect 58494 79662 58546 79714
rect 62750 79662 62802 79714
rect 63086 79662 63138 79714
rect 66446 79662 66498 79714
rect 67454 79662 67506 79714
rect 74174 79662 74226 79714
rect 80334 79662 80386 79714
rect 80670 79662 80722 79714
rect 82126 79662 82178 79714
rect 85262 79662 85314 79714
rect 86270 79662 86322 79714
rect 94558 79662 94610 79714
rect 94894 79662 94946 79714
rect 95790 79662 95842 79714
rect 96126 79662 96178 79714
rect 49534 79550 49586 79602
rect 54686 79550 54738 79602
rect 57934 79550 57986 79602
rect 58270 79550 58322 79602
rect 59054 79550 59106 79602
rect 59502 79550 59554 79602
rect 60510 79550 60562 79602
rect 63310 79550 63362 79602
rect 66782 79550 66834 79602
rect 67230 79550 67282 79602
rect 68126 79550 68178 79602
rect 68686 79550 68738 79602
rect 69582 79550 69634 79602
rect 70478 79550 70530 79602
rect 71598 79550 71650 79602
rect 72494 79550 72546 79602
rect 73502 79550 73554 79602
rect 81454 79550 81506 79602
rect 85598 79550 85650 79602
rect 86046 79550 86098 79602
rect 86830 79550 86882 79602
rect 87502 79550 87554 79602
rect 88398 79550 88450 79602
rect 93326 79550 93378 79602
rect 97582 79550 97634 79602
rect 52446 79438 52498 79490
rect 61182 79438 61234 79490
rect 61630 79438 61682 79490
rect 76302 79438 76354 79490
rect 76750 79438 76802 79490
rect 77198 79438 77250 79490
rect 84254 79438 84306 79490
rect 90414 79438 90466 79490
rect 92542 79438 92594 79490
rect 84478 79326 84530 79378
rect 85038 79326 85090 79378
rect 93998 79326 94050 79378
rect 94334 79326 94386 79378
rect 4478 79158 4530 79210
rect 4582 79158 4634 79210
rect 4686 79158 4738 79210
rect 35198 79158 35250 79210
rect 35302 79158 35354 79210
rect 35406 79158 35458 79210
rect 65918 79158 65970 79210
rect 66022 79158 66074 79210
rect 66126 79158 66178 79210
rect 96638 79158 96690 79210
rect 96742 79158 96794 79210
rect 96846 79158 96898 79210
rect 54574 78878 54626 78930
rect 57374 78878 57426 78930
rect 67230 78878 67282 78930
rect 73838 78878 73890 78930
rect 80446 78878 80498 78930
rect 85262 78878 85314 78930
rect 88958 78878 89010 78930
rect 95678 78878 95730 78930
rect 97806 78878 97858 78930
rect 52110 78766 52162 78818
rect 52446 78766 52498 78818
rect 53342 78766 53394 78818
rect 57822 78766 57874 78818
rect 58270 78766 58322 78818
rect 59390 78766 59442 78818
rect 60398 78766 60450 78818
rect 62302 78766 62354 78818
rect 64318 78766 64370 78818
rect 68574 78766 68626 78818
rect 69582 78766 69634 78818
rect 75966 78766 76018 78818
rect 82014 78766 82066 78818
rect 83022 78766 83074 78818
rect 83806 78766 83858 78818
rect 85710 78766 85762 78818
rect 86158 78766 86210 78818
rect 86718 78766 86770 78818
rect 87502 78766 87554 78818
rect 88398 78766 88450 78818
rect 91646 78766 91698 78818
rect 93214 78766 93266 78818
rect 94894 78766 94946 78818
rect 49310 78654 49362 78706
rect 50654 78654 50706 78706
rect 50766 78654 50818 78706
rect 51662 78654 51714 78706
rect 53566 78654 53618 78706
rect 53678 78654 53730 78706
rect 58830 78654 58882 78706
rect 65102 78654 65154 78706
rect 67790 78654 67842 78706
rect 67902 78654 67954 78706
rect 75182 78654 75234 78706
rect 75518 78654 75570 78706
rect 76302 78654 76354 78706
rect 83358 78654 83410 78706
rect 84030 78654 84082 78706
rect 84142 78654 84194 78706
rect 91870 78654 91922 78706
rect 49758 78542 49810 78594
rect 50206 78542 50258 78594
rect 50990 78542 51042 78594
rect 51326 78542 51378 78594
rect 51550 78542 51602 78594
rect 52334 78542 52386 78594
rect 54238 78542 54290 78594
rect 58382 78542 58434 78594
rect 61294 78542 61346 78594
rect 61742 78542 61794 78594
rect 62638 78542 62690 78594
rect 68126 78542 68178 78594
rect 76190 78542 76242 78594
rect 83246 78542 83298 78594
rect 86270 78542 86322 78594
rect 89518 78542 89570 78594
rect 93550 78542 93602 78594
rect 19838 78374 19890 78426
rect 19942 78374 19994 78426
rect 20046 78374 20098 78426
rect 50558 78374 50610 78426
rect 50662 78374 50714 78426
rect 50766 78374 50818 78426
rect 81278 78374 81330 78426
rect 81382 78374 81434 78426
rect 81486 78374 81538 78426
rect 48862 78206 48914 78258
rect 49982 78206 50034 78258
rect 50766 78206 50818 78258
rect 53678 78206 53730 78258
rect 54126 78206 54178 78258
rect 63422 78206 63474 78258
rect 65326 78206 65378 78258
rect 66334 78206 66386 78258
rect 67678 78206 67730 78258
rect 69806 78206 69858 78258
rect 70030 78206 70082 78258
rect 70590 78206 70642 78258
rect 96350 78206 96402 78258
rect 48302 78094 48354 78146
rect 49646 78094 49698 78146
rect 49758 78094 49810 78146
rect 50430 78094 50482 78146
rect 50542 78094 50594 78146
rect 51326 78094 51378 78146
rect 52110 78094 52162 78146
rect 54910 78094 54962 78146
rect 56590 78094 56642 78146
rect 58046 78094 58098 78146
rect 59278 78094 59330 78146
rect 60286 78094 60338 78146
rect 65550 78094 65602 78146
rect 69022 78094 69074 78146
rect 69358 78094 69410 78146
rect 70142 78094 70194 78146
rect 77310 78094 77362 78146
rect 78318 78094 78370 78146
rect 89406 78094 89458 78146
rect 89518 78094 89570 78146
rect 93550 78094 93602 78146
rect 95454 78094 95506 78146
rect 51214 77982 51266 78034
rect 51550 77982 51602 78034
rect 51886 77982 51938 78034
rect 52222 77982 52274 78034
rect 52670 77982 52722 78034
rect 55022 77982 55074 78034
rect 56366 77982 56418 78034
rect 56702 77982 56754 78034
rect 57822 77982 57874 78034
rect 58158 77982 58210 78034
rect 59726 77982 59778 78034
rect 60062 77982 60114 78034
rect 60958 77982 61010 78034
rect 61518 77982 61570 78034
rect 62302 77982 62354 78034
rect 65662 77982 65714 78034
rect 66110 77982 66162 78034
rect 66446 77982 66498 78034
rect 66894 77982 66946 78034
rect 68014 77982 68066 78034
rect 68462 77982 68514 78034
rect 71598 77982 71650 78034
rect 72046 77982 72098 78034
rect 73950 77982 74002 78034
rect 77758 77982 77810 78034
rect 78094 77982 78146 78034
rect 78766 77982 78818 78034
rect 79326 77982 79378 78034
rect 80334 77982 80386 78034
rect 81454 77982 81506 78034
rect 87614 77982 87666 78034
rect 88398 77982 88450 78034
rect 89182 77982 89234 78034
rect 94334 77982 94386 78034
rect 95230 77982 95282 78034
rect 53118 77870 53170 77922
rect 57374 77870 57426 77922
rect 58606 77870 58658 77922
rect 62974 77870 63026 77922
rect 71038 77870 71090 77922
rect 73278 77870 73330 77922
rect 74622 77870 74674 77922
rect 76750 77870 76802 77922
rect 82126 77870 82178 77922
rect 84254 77870 84306 77922
rect 84702 77870 84754 77922
rect 85486 77870 85538 77922
rect 91422 77870 91474 77922
rect 54910 77758 54962 77810
rect 96014 77758 96066 77810
rect 4478 77590 4530 77642
rect 4582 77590 4634 77642
rect 4686 77590 4738 77642
rect 35198 77590 35250 77642
rect 35302 77590 35354 77642
rect 35406 77590 35458 77642
rect 65918 77590 65970 77642
rect 66022 77590 66074 77642
rect 66126 77590 66178 77642
rect 96638 77590 96690 77642
rect 96742 77590 96794 77642
rect 96846 77590 96898 77642
rect 57486 77422 57538 77474
rect 58270 77422 58322 77474
rect 72830 77422 72882 77474
rect 94334 77422 94386 77474
rect 94894 77422 94946 77474
rect 52670 77310 52722 77362
rect 55134 77310 55186 77362
rect 57262 77310 57314 77362
rect 69246 77310 69298 77362
rect 79886 77310 79938 77362
rect 82238 77310 82290 77362
rect 85262 77310 85314 77362
rect 88734 77310 88786 77362
rect 94670 77310 94722 77362
rect 49870 77198 49922 77250
rect 54350 77198 54402 77250
rect 57710 77198 57762 77250
rect 62078 77198 62130 77250
rect 67902 77198 67954 77250
rect 70814 77198 70866 77250
rect 71822 77198 71874 77250
rect 76526 77198 76578 77250
rect 78878 77198 78930 77250
rect 80446 77198 80498 77250
rect 80782 77198 80834 77250
rect 84366 77198 84418 77250
rect 88174 77198 88226 77250
rect 93326 77198 93378 77250
rect 50542 77086 50594 77138
rect 64318 77086 64370 77138
rect 72158 77086 72210 77138
rect 72718 77086 72770 77138
rect 72830 77086 72882 77138
rect 74958 77086 75010 77138
rect 75518 77086 75570 77138
rect 77198 77086 77250 77138
rect 77534 77086 77586 77138
rect 77982 77086 78034 77138
rect 78206 77086 78258 77138
rect 78318 77086 78370 77138
rect 79214 77086 79266 77138
rect 81454 77086 81506 77138
rect 81790 77086 81842 77138
rect 83022 77086 83074 77138
rect 83134 77086 83186 77138
rect 87390 77086 87442 77138
rect 53342 76974 53394 77026
rect 53790 76974 53842 77026
rect 58158 76974 58210 77026
rect 58606 76974 58658 77026
rect 68350 76974 68402 77026
rect 69694 76974 69746 77026
rect 71262 76974 71314 77026
rect 71934 76974 71986 77026
rect 74286 76974 74338 77026
rect 74622 76974 74674 77026
rect 74846 76974 74898 77026
rect 75854 76974 75906 77026
rect 77422 76974 77474 77026
rect 81678 76974 81730 77026
rect 83358 76974 83410 77026
rect 84030 76974 84082 77026
rect 84254 76974 84306 77026
rect 90862 76974 90914 77026
rect 92542 76974 92594 77026
rect 93550 76974 93602 77026
rect 95006 76974 95058 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 81278 76806 81330 76858
rect 81382 76806 81434 76858
rect 81486 76806 81538 76858
rect 58382 76638 58434 76690
rect 58942 76638 58994 76690
rect 63534 76638 63586 76690
rect 64542 76638 64594 76690
rect 65438 76638 65490 76690
rect 67006 76638 67058 76690
rect 76974 76638 77026 76690
rect 77758 76638 77810 76690
rect 78542 76638 78594 76690
rect 80222 76638 80274 76690
rect 87278 76638 87330 76690
rect 87614 76638 87666 76690
rect 57598 76526 57650 76578
rect 57710 76526 57762 76578
rect 64766 76526 64818 76578
rect 66446 76526 66498 76578
rect 66558 76526 66610 76578
rect 67230 76526 67282 76578
rect 74398 76526 74450 76578
rect 81454 76526 81506 76578
rect 82238 76526 82290 76578
rect 82798 76526 82850 76578
rect 84254 76526 84306 76578
rect 87054 76526 87106 76578
rect 90302 76526 90354 76578
rect 52894 76414 52946 76466
rect 58494 76414 58546 76466
rect 64430 76414 64482 76466
rect 65774 76414 65826 76466
rect 67342 76414 67394 76466
rect 68126 76414 68178 76466
rect 71598 76414 71650 76466
rect 73726 76414 73778 76466
rect 81230 76414 81282 76466
rect 81566 76414 81618 76466
rect 82350 76414 82402 76466
rect 83582 76414 83634 76466
rect 86942 76414 86994 76466
rect 90638 76414 90690 76466
rect 91870 76414 91922 76466
rect 50878 76302 50930 76354
rect 56478 76302 56530 76354
rect 63870 76302 63922 76354
rect 68910 76302 68962 76354
rect 71038 76302 71090 76354
rect 72158 76302 72210 76354
rect 72606 76302 72658 76354
rect 76526 76302 76578 76354
rect 80558 76302 80610 76354
rect 86382 76302 86434 76354
rect 94894 76302 94946 76354
rect 97134 76302 97186 76354
rect 57598 76190 57650 76242
rect 58382 76190 58434 76242
rect 66446 76190 66498 76242
rect 82238 76190 82290 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 96638 76022 96690 76074
rect 96742 76022 96794 76074
rect 96846 76022 96898 76074
rect 67566 75854 67618 75906
rect 68126 75854 68178 75906
rect 97134 75854 97186 75906
rect 50542 75742 50594 75794
rect 52670 75742 52722 75794
rect 56702 75742 56754 75794
rect 58046 75742 58098 75794
rect 60174 75742 60226 75794
rect 62974 75742 63026 75794
rect 64542 75742 64594 75794
rect 66670 75742 66722 75794
rect 67566 75742 67618 75794
rect 70142 75742 70194 75794
rect 70590 75742 70642 75794
rect 71262 75742 71314 75794
rect 73390 75742 73442 75794
rect 73726 75742 73778 75794
rect 79774 75742 79826 75794
rect 81902 75742 81954 75794
rect 86718 75742 86770 75794
rect 90302 75742 90354 75794
rect 92430 75742 92482 75794
rect 93214 75742 93266 75794
rect 95342 75742 95394 75794
rect 49870 75630 49922 75682
rect 53790 75630 53842 75682
rect 57374 75630 57426 75682
rect 63758 75630 63810 75682
rect 67118 75630 67170 75682
rect 68014 75630 68066 75682
rect 74622 75630 74674 75682
rect 76302 75630 76354 75682
rect 79102 75630 79154 75682
rect 82350 75630 82402 75682
rect 82686 75630 82738 75682
rect 83470 75630 83522 75682
rect 84590 75630 84642 75682
rect 85598 75630 85650 75682
rect 86046 75630 86098 75682
rect 86382 75630 86434 75682
rect 89518 75630 89570 75682
rect 96014 75630 96066 75682
rect 54574 75518 54626 75570
rect 62526 75518 62578 75570
rect 69358 75518 69410 75570
rect 69694 75518 69746 75570
rect 74286 75518 74338 75570
rect 75070 75518 75122 75570
rect 75406 75518 75458 75570
rect 75966 75518 76018 75570
rect 76078 75518 76130 75570
rect 84254 75518 84306 75570
rect 85262 75518 85314 75570
rect 85374 75518 85426 75570
rect 86158 75518 86210 75570
rect 97358 75518 97410 75570
rect 97806 75518 97858 75570
rect 62190 75406 62242 75458
rect 74398 75406 74450 75458
rect 82574 75406 82626 75458
rect 83134 75406 83186 75458
rect 83358 75406 83410 75458
rect 84366 75406 84418 75458
rect 89070 75406 89122 75458
rect 96798 75406 96850 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 81278 75238 81330 75290
rect 81382 75238 81434 75290
rect 81486 75238 81538 75290
rect 53342 75070 53394 75122
rect 53566 75070 53618 75122
rect 54126 75070 54178 75122
rect 54910 75070 54962 75122
rect 55134 75070 55186 75122
rect 55694 75070 55746 75122
rect 57374 75070 57426 75122
rect 57822 75070 57874 75122
rect 65438 75070 65490 75122
rect 66222 75070 66274 75122
rect 70590 75070 70642 75122
rect 74622 75070 74674 75122
rect 76078 75070 76130 75122
rect 85150 75070 85202 75122
rect 91422 75070 91474 75122
rect 93438 75070 93490 75122
rect 50766 74958 50818 75010
rect 54350 74958 54402 75010
rect 55918 74958 55970 75010
rect 56030 74958 56082 75010
rect 65774 74958 65826 75010
rect 71486 74958 71538 75010
rect 75070 74958 75122 75010
rect 88510 74958 88562 75010
rect 89966 74958 90018 75010
rect 90526 74958 90578 75010
rect 91982 74958 92034 75010
rect 92318 74958 92370 75010
rect 93998 74958 94050 75010
rect 94334 74958 94386 75010
rect 95566 74958 95618 75010
rect 95902 74958 95954 75010
rect 49982 74846 50034 74898
rect 53678 74846 53730 74898
rect 54462 74846 54514 74898
rect 55246 74846 55298 74898
rect 60622 74846 60674 74898
rect 64318 74846 64370 74898
rect 67006 74846 67058 74898
rect 70926 74846 70978 74898
rect 71710 74846 71762 74898
rect 74286 74846 74338 74898
rect 81790 74846 81842 74898
rect 88286 74846 88338 74898
rect 89406 74846 89458 74898
rect 52894 74734 52946 74786
rect 56478 74734 56530 74786
rect 61294 74734 61346 74786
rect 63422 74734 63474 74786
rect 63982 74734 64034 74786
rect 67790 74734 67842 74786
rect 69918 74734 69970 74786
rect 72270 74734 72322 74786
rect 73726 74734 73778 74786
rect 75742 74734 75794 74786
rect 81342 74734 81394 74786
rect 82574 74734 82626 74786
rect 84702 74734 84754 74786
rect 89742 74734 89794 74786
rect 96350 74734 96402 74786
rect 97134 74734 97186 74786
rect 91758 74622 91810 74674
rect 93774 74622 93826 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 96638 74454 96690 74506
rect 96742 74454 96794 74506
rect 96846 74454 96898 74506
rect 82574 74286 82626 74338
rect 82910 74286 82962 74338
rect 50206 74174 50258 74226
rect 53342 74174 53394 74226
rect 53902 74174 53954 74226
rect 54350 74174 54402 74226
rect 54798 74174 54850 74226
rect 67566 74174 67618 74226
rect 82238 74174 82290 74226
rect 82686 74174 82738 74226
rect 84366 74174 84418 74226
rect 88622 74174 88674 74226
rect 90750 74174 90802 74226
rect 91646 74174 91698 74226
rect 92094 74174 92146 74226
rect 93102 74174 93154 74226
rect 93550 74174 93602 74226
rect 95678 74174 95730 74226
rect 97806 74174 97858 74226
rect 50654 74062 50706 74114
rect 51326 74062 51378 74114
rect 51662 74062 51714 74114
rect 52110 74062 52162 74114
rect 52446 74062 52498 74114
rect 60398 74062 60450 74114
rect 61518 74062 61570 74114
rect 61854 74062 61906 74114
rect 62414 74062 62466 74114
rect 63870 74062 63922 74114
rect 69806 74062 69858 74114
rect 74846 74062 74898 74114
rect 76078 74062 76130 74114
rect 76526 74062 76578 74114
rect 83022 74062 83074 74114
rect 83358 74062 83410 74114
rect 87838 74062 87890 74114
rect 94894 74062 94946 74114
rect 50990 73950 51042 74002
rect 59726 73950 59778 74002
rect 60622 73950 60674 74002
rect 62638 73950 62690 74002
rect 69470 73950 69522 74002
rect 70030 73950 70082 74002
rect 70590 73950 70642 74002
rect 71934 73950 71986 74002
rect 72270 73950 72322 74002
rect 72718 73950 72770 74002
rect 77422 73950 77474 74002
rect 78542 73950 78594 74002
rect 83806 73950 83858 74002
rect 91310 73950 91362 74002
rect 50766 73838 50818 73890
rect 51550 73838 51602 73890
rect 52334 73838 52386 73890
rect 71262 73838 71314 73890
rect 75070 73838 75122 73890
rect 78206 73838 78258 73890
rect 83246 73838 83298 73890
rect 93998 73838 94050 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 81278 73670 81330 73722
rect 81382 73670 81434 73722
rect 81486 73670 81538 73722
rect 58270 73502 58322 73554
rect 59502 73502 59554 73554
rect 65326 73502 65378 73554
rect 68238 73502 68290 73554
rect 79326 73502 79378 73554
rect 91086 73502 91138 73554
rect 56030 73390 56082 73442
rect 62190 73390 62242 73442
rect 68574 73390 68626 73442
rect 75070 73390 75122 73442
rect 78318 73390 78370 73442
rect 78766 73390 78818 73442
rect 81790 73390 81842 73442
rect 83246 73390 83298 73442
rect 88174 73390 88226 73442
rect 89966 73390 90018 73442
rect 90526 73390 90578 73442
rect 91982 73390 92034 73442
rect 93662 73390 93714 73442
rect 95790 73390 95842 73442
rect 96350 73390 96402 73442
rect 97246 73390 97298 73442
rect 56366 73278 56418 73330
rect 61518 73278 61570 73330
rect 73726 73278 73778 73330
rect 74398 73278 74450 73330
rect 81566 73278 81618 73330
rect 83022 73278 83074 73330
rect 88510 73278 88562 73330
rect 89406 73278 89458 73330
rect 91758 73278 91810 73330
rect 95230 73278 95282 73330
rect 97582 73278 97634 73330
rect 51326 73166 51378 73218
rect 51886 73166 51938 73218
rect 57486 73166 57538 73218
rect 57822 73166 57874 73218
rect 60846 73166 60898 73218
rect 64318 73166 64370 73218
rect 71150 73166 71202 73218
rect 72494 73166 72546 73218
rect 73390 73166 73442 73218
rect 77198 73166 77250 73218
rect 79998 73166 80050 73218
rect 94222 73166 94274 73218
rect 94670 73166 94722 73218
rect 78990 73054 79042 73106
rect 89742 73054 89794 73106
rect 94222 73054 94274 73106
rect 94894 73054 94946 73106
rect 95566 73054 95618 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 96638 72886 96690 72938
rect 96742 72886 96794 72938
rect 96846 72886 96898 72938
rect 58046 72718 58098 72770
rect 62078 72718 62130 72770
rect 64766 72718 64818 72770
rect 74846 72718 74898 72770
rect 59726 72606 59778 72658
rect 71710 72606 71762 72658
rect 73502 72606 73554 72658
rect 77870 72606 77922 72658
rect 94894 72606 94946 72658
rect 97022 72606 97074 72658
rect 49758 72494 49810 72546
rect 56478 72494 56530 72546
rect 57150 72494 57202 72546
rect 58382 72494 58434 72546
rect 59166 72494 59218 72546
rect 60398 72494 60450 72546
rect 61742 72494 61794 72546
rect 62750 72494 62802 72546
rect 64430 72494 64482 72546
rect 72270 72494 72322 72546
rect 73950 72494 74002 72546
rect 75182 72494 75234 72546
rect 75630 72494 75682 72546
rect 83918 72494 83970 72546
rect 87166 72494 87218 72546
rect 97694 72494 97746 72546
rect 55470 72382 55522 72434
rect 56142 72382 56194 72434
rect 57262 72382 57314 72434
rect 59054 72382 59106 72434
rect 62862 72382 62914 72434
rect 63646 72382 63698 72434
rect 64206 72382 64258 72434
rect 70814 72382 70866 72434
rect 75966 72382 76018 72434
rect 78990 72382 79042 72434
rect 89182 72382 89234 72434
rect 49982 72270 50034 72322
rect 54686 72270 54738 72322
rect 55134 72270 55186 72322
rect 60622 72270 60674 72322
rect 65326 72270 65378 72322
rect 65774 72270 65826 72322
rect 69246 72270 69298 72322
rect 70478 72270 70530 72322
rect 72830 72270 72882 72322
rect 76526 72270 76578 72322
rect 77198 72270 77250 72322
rect 84478 72270 84530 72322
rect 86606 72270 86658 72322
rect 94110 72270 94162 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 81278 72102 81330 72154
rect 81382 72102 81434 72154
rect 81486 72102 81538 72154
rect 50430 71934 50482 71986
rect 63646 71934 63698 71986
rect 73838 71934 73890 71986
rect 51550 71822 51602 71874
rect 54574 71822 54626 71874
rect 68910 71822 68962 71874
rect 70254 71822 70306 71874
rect 78430 71822 78482 71874
rect 82126 71822 82178 71874
rect 92542 71822 92594 71874
rect 51438 71710 51490 71762
rect 53790 71710 53842 71762
rect 62750 71710 62802 71762
rect 68686 71710 68738 71762
rect 69582 71710 69634 71762
rect 77646 71710 77698 71762
rect 81342 71710 81394 71762
rect 89854 71710 89906 71762
rect 52110 71598 52162 71650
rect 52670 71598 52722 71650
rect 53342 71598 53394 71650
rect 56702 71598 56754 71650
rect 58830 71598 58882 71650
rect 63198 71598 63250 71650
rect 66110 71598 66162 71650
rect 68014 71598 68066 71650
rect 72382 71598 72434 71650
rect 73278 71598 73330 71650
rect 74286 71598 74338 71650
rect 74846 71598 74898 71650
rect 75294 71598 75346 71650
rect 75742 71598 75794 71650
rect 76302 71598 76354 71650
rect 76638 71598 76690 71650
rect 80558 71598 80610 71650
rect 84254 71598 84306 71650
rect 95566 71598 95618 71650
rect 50766 71486 50818 71538
rect 74846 71486 74898 71538
rect 75294 71486 75346 71538
rect 76750 71486 76802 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 96638 71318 96690 71370
rect 96742 71318 96794 71370
rect 96846 71318 96898 71370
rect 82014 71150 82066 71202
rect 82350 71150 82402 71202
rect 85374 71150 85426 71202
rect 85710 71150 85762 71202
rect 92318 71150 92370 71202
rect 51662 71038 51714 71090
rect 55806 71038 55858 71090
rect 57934 71038 57986 71090
rect 62190 71038 62242 71090
rect 64318 71038 64370 71090
rect 67230 71038 67282 71090
rect 71374 71038 71426 71090
rect 77198 71038 77250 71090
rect 80334 71038 80386 71090
rect 80782 71038 80834 71090
rect 88398 71038 88450 71090
rect 90526 71038 90578 71090
rect 93662 71038 93714 71090
rect 93998 71038 94050 71090
rect 96462 71038 96514 71090
rect 48862 70926 48914 70978
rect 55134 70926 55186 70978
rect 58942 70926 58994 70978
rect 61518 70926 61570 70978
rect 69358 70926 69410 70978
rect 75294 70926 75346 70978
rect 76078 70926 76130 70978
rect 83022 70926 83074 70978
rect 87726 70926 87778 70978
rect 91310 70926 91362 70978
rect 91982 70926 92034 70978
rect 93102 70926 93154 70978
rect 47854 70814 47906 70866
rect 48190 70814 48242 70866
rect 49534 70814 49586 70866
rect 53566 70814 53618 70866
rect 53902 70814 53954 70866
rect 59166 70814 59218 70866
rect 59502 70814 59554 70866
rect 65662 70814 65714 70866
rect 66334 70814 66386 70866
rect 66670 70814 66722 70866
rect 68238 70814 68290 70866
rect 68574 70814 68626 70866
rect 82910 70814 82962 70866
rect 85934 70814 85986 70866
rect 86270 70814 86322 70866
rect 91198 70814 91250 70866
rect 94782 70814 94834 70866
rect 95118 70814 95170 70866
rect 95678 70814 95730 70866
rect 52110 70702 52162 70754
rect 52670 70702 52722 70754
rect 58606 70702 58658 70754
rect 60286 70702 60338 70754
rect 64766 70702 64818 70754
rect 65326 70702 65378 70754
rect 67790 70702 67842 70754
rect 75518 70702 75570 70754
rect 76414 70702 76466 70754
rect 77758 70702 77810 70754
rect 81454 70702 81506 70754
rect 83694 70702 83746 70754
rect 84590 70702 84642 70754
rect 87054 70702 87106 70754
rect 96014 70702 96066 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 81278 70534 81330 70586
rect 81382 70534 81434 70586
rect 81486 70534 81538 70586
rect 63870 70366 63922 70418
rect 66222 70366 66274 70418
rect 71486 70366 71538 70418
rect 72606 70366 72658 70418
rect 81230 70366 81282 70418
rect 88062 70366 88114 70418
rect 89294 70366 89346 70418
rect 94782 70366 94834 70418
rect 56478 70254 56530 70306
rect 58494 70254 58546 70306
rect 66782 70254 66834 70306
rect 67342 70254 67394 70306
rect 68910 70254 68962 70306
rect 76190 70254 76242 70306
rect 83246 70254 83298 70306
rect 90302 70254 90354 70306
rect 93102 70254 93154 70306
rect 95342 70254 95394 70306
rect 95678 70254 95730 70306
rect 52894 70142 52946 70194
rect 58718 70142 58770 70194
rect 59278 70142 59330 70194
rect 60622 70142 60674 70194
rect 68126 70142 68178 70194
rect 72046 70142 72098 70194
rect 76974 70142 77026 70194
rect 77646 70142 77698 70194
rect 82574 70142 82626 70194
rect 87166 70142 87218 70194
rect 89630 70142 89682 70194
rect 90190 70142 90242 70194
rect 90526 70142 90578 70194
rect 93886 70142 93938 70194
rect 96462 70142 96514 70194
rect 59726 70030 59778 70082
rect 61294 70030 61346 70082
rect 63422 70030 63474 70082
rect 71038 70030 71090 70082
rect 73390 70030 73442 70082
rect 74062 70030 74114 70082
rect 78318 70030 78370 70082
rect 80446 70030 80498 70082
rect 85374 70030 85426 70082
rect 87726 70030 87778 70082
rect 88510 70030 88562 70082
rect 90974 70030 91026 70082
rect 95118 70030 95170 70082
rect 97134 70030 97186 70082
rect 57598 69918 57650 69970
rect 57934 69918 57986 69970
rect 59054 69918 59106 69970
rect 59838 69918 59890 69970
rect 66558 69918 66610 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 96638 69750 96690 69802
rect 96742 69750 96794 69802
rect 96846 69750 96898 69802
rect 70254 69582 70306 69634
rect 72158 69582 72210 69634
rect 72494 69582 72546 69634
rect 75742 69582 75794 69634
rect 84366 69582 84418 69634
rect 52446 69470 52498 69522
rect 56478 69470 56530 69522
rect 59950 69470 60002 69522
rect 60398 69470 60450 69522
rect 63870 69470 63922 69522
rect 69246 69470 69298 69522
rect 81230 69470 81282 69522
rect 82686 69470 82738 69522
rect 86046 69470 86098 69522
rect 88174 69470 88226 69522
rect 89518 69470 89570 69522
rect 94110 69470 94162 69522
rect 94894 69470 94946 69522
rect 97022 69470 97074 69522
rect 49534 69358 49586 69410
rect 53678 69358 53730 69410
rect 57150 69358 57202 69410
rect 65438 69358 65490 69410
rect 70590 69358 70642 69410
rect 71262 69358 71314 69410
rect 73278 69358 73330 69410
rect 75406 69358 75458 69410
rect 78206 69358 78258 69410
rect 79102 69358 79154 69410
rect 81902 69358 81954 69410
rect 84478 69358 84530 69410
rect 85262 69358 85314 69410
rect 89070 69358 89122 69410
rect 92430 69358 92482 69410
rect 93438 69358 93490 69410
rect 97694 69358 97746 69410
rect 50318 69246 50370 69298
rect 54350 69246 54402 69298
rect 57822 69246 57874 69298
rect 67566 69246 67618 69298
rect 67678 69246 67730 69298
rect 68574 69246 68626 69298
rect 71374 69246 71426 69298
rect 73054 69246 73106 69298
rect 74846 69246 74898 69298
rect 75182 69246 75234 69298
rect 77422 69246 77474 69298
rect 77982 69246 78034 69298
rect 82126 69246 82178 69298
rect 83246 69246 83298 69298
rect 83358 69246 83410 69298
rect 88734 69246 88786 69298
rect 88846 69246 88898 69298
rect 91646 69246 91698 69298
rect 93214 69246 93266 69298
rect 67902 69134 67954 69186
rect 68238 69134 68290 69186
rect 68462 69134 68514 69186
rect 73950 69134 74002 69186
rect 76302 69134 76354 69186
rect 78542 69134 78594 69186
rect 79550 69134 79602 69186
rect 79998 69134 80050 69186
rect 83582 69134 83634 69186
rect 84366 69134 84418 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 81278 68966 81330 69018
rect 81382 68966 81434 69018
rect 81486 68966 81538 69018
rect 50206 68798 50258 68850
rect 52670 68798 52722 68850
rect 53678 68798 53730 68850
rect 54238 68798 54290 68850
rect 55134 68798 55186 68850
rect 56478 68798 56530 68850
rect 57374 68798 57426 68850
rect 60622 68798 60674 68850
rect 61182 68798 61234 68850
rect 65550 68798 65602 68850
rect 73726 68798 73778 68850
rect 74846 68798 74898 68850
rect 77198 68798 77250 68850
rect 90526 68798 90578 68850
rect 51326 68686 51378 68738
rect 52110 68686 52162 68738
rect 54574 68686 54626 68738
rect 63310 68686 63362 68738
rect 75742 68686 75794 68738
rect 78094 68686 78146 68738
rect 79214 68686 79266 68738
rect 79998 68686 80050 68738
rect 89630 68686 89682 68738
rect 96238 68686 96290 68738
rect 51214 68574 51266 68626
rect 51886 68574 51938 68626
rect 52222 68574 52274 68626
rect 55358 68574 55410 68626
rect 56254 68574 56306 68626
rect 61518 68574 61570 68626
rect 62190 68574 62242 68626
rect 63198 68574 63250 68626
rect 63870 68574 63922 68626
rect 66110 68574 66162 68626
rect 74286 68574 74338 68626
rect 75182 68574 75234 68626
rect 76302 68574 76354 68626
rect 76974 68574 77026 68626
rect 77758 68574 77810 68626
rect 79102 68574 79154 68626
rect 79438 68574 79490 68626
rect 79886 68574 79938 68626
rect 87390 68574 87442 68626
rect 89406 68574 89458 68626
rect 90190 68574 90242 68626
rect 91198 68574 91250 68626
rect 53118 68462 53170 68514
rect 64318 68462 64370 68514
rect 66894 68462 66946 68514
rect 69022 68462 69074 68514
rect 69582 68462 69634 68514
rect 69918 68462 69970 68514
rect 70590 68462 70642 68514
rect 71038 68462 71090 68514
rect 71374 68462 71426 68514
rect 71934 68462 71986 68514
rect 72494 68462 72546 68514
rect 78654 68462 78706 68514
rect 83470 68462 83522 68514
rect 50542 68350 50594 68402
rect 52446 68350 52498 68402
rect 53006 68350 53058 68402
rect 62526 68350 62578 68402
rect 79998 68350 80050 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 96638 68182 96690 68234
rect 96742 68182 96794 68234
rect 96846 68182 96898 68234
rect 52110 68014 52162 68066
rect 52558 68014 52610 68066
rect 61854 68014 61906 68066
rect 68462 68014 68514 68066
rect 49646 67902 49698 67954
rect 51774 67902 51826 67954
rect 59390 67902 59442 67954
rect 63198 67902 63250 67954
rect 64878 67902 64930 67954
rect 67006 67902 67058 67954
rect 69246 67902 69298 67954
rect 72606 67902 72658 67954
rect 73390 67902 73442 67954
rect 75742 67902 75794 67954
rect 76190 67902 76242 67954
rect 77534 67902 77586 67954
rect 88174 67902 88226 67954
rect 88734 67902 88786 67954
rect 90862 67902 90914 67954
rect 92094 67902 92146 67954
rect 93550 67902 93602 67954
rect 95678 67902 95730 67954
rect 48974 67790 49026 67842
rect 62302 67790 62354 67842
rect 64094 67790 64146 67842
rect 67454 67790 67506 67842
rect 67790 67790 67842 67842
rect 72494 67790 72546 67842
rect 73838 67790 73890 67842
rect 82574 67790 82626 67842
rect 83022 67790 83074 67842
rect 84254 67790 84306 67842
rect 85262 67790 85314 67842
rect 91534 67790 91586 67842
rect 96350 67790 96402 67842
rect 97358 67790 97410 67842
rect 60622 67678 60674 67730
rect 61518 67678 61570 67730
rect 62638 67678 62690 67730
rect 67678 67678 67730 67730
rect 68462 67678 68514 67730
rect 68574 67678 68626 67730
rect 72830 67678 72882 67730
rect 83582 67678 83634 67730
rect 83694 67678 83746 67730
rect 86046 67678 86098 67730
rect 52222 67566 52274 67618
rect 52670 67566 52722 67618
rect 53342 67566 53394 67618
rect 53790 67566 53842 67618
rect 54798 67566 54850 67618
rect 60286 67566 60338 67618
rect 69918 67566 69970 67618
rect 70590 67566 70642 67618
rect 71150 67566 71202 67618
rect 71598 67566 71650 67618
rect 72046 67566 72098 67618
rect 74510 67566 74562 67618
rect 74958 67566 75010 67618
rect 75406 67566 75458 67618
rect 83918 67566 83970 67618
rect 96910 67566 96962 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 81278 67398 81330 67450
rect 81382 67398 81434 67450
rect 81486 67398 81538 67450
rect 50318 67230 50370 67282
rect 51998 67230 52050 67282
rect 52558 67230 52610 67282
rect 52782 67230 52834 67282
rect 63534 67230 63586 67282
rect 71822 67230 71874 67282
rect 73390 67230 73442 67282
rect 74510 67230 74562 67282
rect 76078 67230 76130 67282
rect 83806 67230 83858 67282
rect 85374 67230 85426 67282
rect 86494 67230 86546 67282
rect 49758 67118 49810 67170
rect 51102 67118 51154 67170
rect 51214 67118 51266 67170
rect 51886 67118 51938 67170
rect 52894 67118 52946 67170
rect 53790 67118 53842 67170
rect 54238 67118 54290 67170
rect 60510 67118 60562 67170
rect 63086 67118 63138 67170
rect 67342 67118 67394 67170
rect 69918 67118 69970 67170
rect 70142 67118 70194 67170
rect 70254 67118 70306 67170
rect 73950 67118 74002 67170
rect 75966 67118 76018 67170
rect 77086 67118 77138 67170
rect 81230 67118 81282 67170
rect 81454 67118 81506 67170
rect 83246 67118 83298 67170
rect 84254 67118 84306 67170
rect 84702 67118 84754 67170
rect 85150 67118 85202 67170
rect 85486 67118 85538 67170
rect 86718 67118 86770 67170
rect 87726 67118 87778 67170
rect 91534 67118 91586 67170
rect 95342 67118 95394 67170
rect 96350 67118 96402 67170
rect 48862 67006 48914 67058
rect 50094 67006 50146 67058
rect 50430 67006 50482 67058
rect 51438 67006 51490 67058
rect 52222 67006 52274 67058
rect 59838 67006 59890 67058
rect 66558 67006 66610 67058
rect 72158 67006 72210 67058
rect 74734 67006 74786 67058
rect 76750 67006 76802 67058
rect 77646 67006 77698 67058
rect 81566 67006 81618 67058
rect 83134 67006 83186 67058
rect 86382 67006 86434 67058
rect 87838 67006 87890 67058
rect 93998 67006 94050 67058
rect 95230 67006 95282 67058
rect 48302 66894 48354 66946
rect 53454 66894 53506 66946
rect 58718 66894 58770 66946
rect 59054 66894 59106 66946
rect 62638 66894 62690 66946
rect 69470 66894 69522 66946
rect 70702 66894 70754 66946
rect 71150 66894 71202 66946
rect 72718 66894 72770 66946
rect 75406 66894 75458 66946
rect 78430 66894 78482 66946
rect 80558 66894 80610 66946
rect 82014 66894 82066 66946
rect 87054 66894 87106 66946
rect 88286 66894 88338 66946
rect 96014 66894 96066 66946
rect 97134 66894 97186 66946
rect 97582 66894 97634 66946
rect 73726 66782 73778 66834
rect 76078 66782 76130 66834
rect 83246 66782 83298 66834
rect 87726 66782 87778 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 96638 66614 96690 66666
rect 96742 66614 96794 66666
rect 96846 66614 96898 66666
rect 65998 66446 66050 66498
rect 74062 66446 74114 66498
rect 90862 66446 90914 66498
rect 56478 66334 56530 66386
rect 57038 66334 57090 66386
rect 58270 66334 58322 66386
rect 63310 66334 63362 66386
rect 67790 66334 67842 66386
rect 73054 66334 73106 66386
rect 79326 66334 79378 66386
rect 81454 66334 81506 66386
rect 81902 66334 81954 66386
rect 82350 66334 82402 66386
rect 85150 66334 85202 66386
rect 88062 66334 88114 66386
rect 90190 66334 90242 66386
rect 91870 66334 91922 66386
rect 94110 66334 94162 66386
rect 97582 66334 97634 66386
rect 98030 66334 98082 66386
rect 49534 66222 49586 66274
rect 52558 66222 52610 66274
rect 53566 66222 53618 66274
rect 58942 66222 58994 66274
rect 60398 66222 60450 66274
rect 61630 66222 61682 66274
rect 61966 66222 62018 66274
rect 66558 66222 66610 66274
rect 67566 66222 67618 66274
rect 68574 66222 68626 66274
rect 69358 66222 69410 66274
rect 74062 66222 74114 66274
rect 75518 66222 75570 66274
rect 77422 66222 77474 66274
rect 78542 66222 78594 66274
rect 85822 66222 85874 66274
rect 87390 66222 87442 66274
rect 94670 66222 94722 66274
rect 49198 66110 49250 66162
rect 50094 66110 50146 66162
rect 50206 66110 50258 66162
rect 50990 66110 51042 66162
rect 51662 66110 51714 66162
rect 51774 66110 51826 66162
rect 54350 66110 54402 66162
rect 58830 66110 58882 66162
rect 62302 66110 62354 66162
rect 62638 66110 62690 66162
rect 66782 66110 66834 66162
rect 67902 66110 67954 66162
rect 69694 66110 69746 66162
rect 73726 66110 73778 66162
rect 74622 66110 74674 66162
rect 74958 66110 75010 66162
rect 75854 66110 75906 66162
rect 84254 66110 84306 66162
rect 84366 66110 84418 66162
rect 90974 66110 91026 66162
rect 91422 66110 91474 66162
rect 93214 66110 93266 66162
rect 93550 66110 93602 66162
rect 95454 66110 95506 66162
rect 49310 65998 49362 66050
rect 49870 65998 49922 66050
rect 50654 65998 50706 66050
rect 50878 65998 50930 66050
rect 51438 65998 51490 66050
rect 52222 65998 52274 66050
rect 52446 65998 52498 66050
rect 58606 65998 58658 66050
rect 59502 65998 59554 66050
rect 60622 65998 60674 66050
rect 64990 65998 65042 66050
rect 65662 65998 65714 66050
rect 67678 65998 67730 66050
rect 68014 65998 68066 66050
rect 69470 65998 69522 66050
rect 70478 65998 70530 66050
rect 70926 65998 70978 66050
rect 71262 65998 71314 66050
rect 71710 65998 71762 66050
rect 72606 65998 72658 66050
rect 76302 65998 76354 66050
rect 77646 65998 77698 66050
rect 82798 65998 82850 66050
rect 83582 65998 83634 66050
rect 84030 65998 84082 66050
rect 85934 65998 85986 66050
rect 86158 65998 86210 66050
rect 86494 65998 86546 66050
rect 90862 65998 90914 66050
rect 92542 65998 92594 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 81278 65830 81330 65882
rect 81382 65830 81434 65882
rect 81486 65830 81538 65882
rect 53790 65662 53842 65714
rect 54014 65662 54066 65714
rect 55246 65662 55298 65714
rect 63310 65662 63362 65714
rect 73502 65662 73554 65714
rect 79102 65662 79154 65714
rect 79774 65662 79826 65714
rect 88062 65662 88114 65714
rect 90190 65662 90242 65714
rect 90862 65662 90914 65714
rect 91310 65662 91362 65714
rect 94558 65662 94610 65714
rect 50318 65550 50370 65602
rect 53118 65550 53170 65602
rect 53230 65550 53282 65602
rect 54126 65550 54178 65602
rect 55022 65550 55074 65602
rect 58606 65550 58658 65602
rect 58718 65550 58770 65602
rect 60734 65550 60786 65602
rect 64318 65550 64370 65602
rect 64654 65550 64706 65602
rect 66334 65550 66386 65602
rect 73950 65550 74002 65602
rect 75966 65550 76018 65602
rect 77758 65550 77810 65602
rect 79662 65550 79714 65602
rect 86718 65550 86770 65602
rect 86830 65550 86882 65602
rect 89406 65550 89458 65602
rect 89518 65550 89570 65602
rect 90302 65550 90354 65602
rect 96350 65550 96402 65602
rect 49646 65438 49698 65490
rect 54574 65438 54626 65490
rect 55358 65438 55410 65490
rect 55806 65438 55858 65490
rect 57598 65438 57650 65490
rect 57822 65438 57874 65490
rect 58158 65438 58210 65490
rect 58942 65438 58994 65490
rect 59950 65438 60002 65490
rect 69246 65438 69298 65490
rect 71150 65438 71202 65490
rect 71598 65438 71650 65490
rect 74958 65438 75010 65490
rect 77198 65438 77250 65490
rect 78094 65438 78146 65490
rect 78878 65438 78930 65490
rect 79998 65438 80050 65490
rect 83246 65438 83298 65490
rect 83918 65438 83970 65490
rect 88174 65438 88226 65490
rect 89182 65438 89234 65490
rect 89966 65438 90018 65490
rect 94334 65438 94386 65490
rect 96126 65438 96178 65490
rect 52446 65326 52498 65378
rect 56702 65326 56754 65378
rect 57934 65326 57986 65378
rect 59278 65326 59330 65378
rect 62862 65326 62914 65378
rect 72046 65326 72098 65378
rect 72718 65326 72770 65378
rect 80334 65326 80386 65378
rect 81230 65326 81282 65378
rect 81790 65326 81842 65378
rect 82238 65326 82290 65378
rect 82686 65326 82738 65378
rect 86046 65326 86098 65378
rect 87390 65326 87442 65378
rect 93774 65326 93826 65378
rect 53118 65214 53170 65266
rect 70926 65214 70978 65266
rect 71486 65214 71538 65266
rect 71710 65214 71762 65266
rect 71934 65214 71986 65266
rect 86718 65214 86770 65266
rect 88062 65214 88114 65266
rect 95230 65214 95282 65266
rect 95566 65214 95618 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 96638 65046 96690 65098
rect 96742 65046 96794 65098
rect 96846 65046 96898 65098
rect 81566 64878 81618 64930
rect 82238 64878 82290 64930
rect 49534 64766 49586 64818
rect 51662 64766 51714 64818
rect 54126 64766 54178 64818
rect 54574 64766 54626 64818
rect 55470 64766 55522 64818
rect 56366 64766 56418 64818
rect 61294 64766 61346 64818
rect 61742 64766 61794 64818
rect 64766 64766 64818 64818
rect 66894 64766 66946 64818
rect 67790 64766 67842 64818
rect 68126 64766 68178 64818
rect 72046 64766 72098 64818
rect 81566 64766 81618 64818
rect 81902 64766 81954 64818
rect 87054 64766 87106 64818
rect 88622 64766 88674 64818
rect 90750 64766 90802 64818
rect 94222 64766 94274 64818
rect 97694 64766 97746 64818
rect 48862 64654 48914 64706
rect 52110 64654 52162 64706
rect 53342 64654 53394 64706
rect 53678 64654 53730 64706
rect 58046 64654 58098 64706
rect 59838 64654 59890 64706
rect 60622 64654 60674 64706
rect 64094 64654 64146 64706
rect 69694 64654 69746 64706
rect 70814 64654 70866 64706
rect 71262 64654 71314 64706
rect 71598 64654 71650 64706
rect 74398 64654 74450 64706
rect 76414 64654 76466 64706
rect 79998 64654 80050 64706
rect 80782 64654 80834 64706
rect 83246 64654 83298 64706
rect 84254 64654 84306 64706
rect 85486 64654 85538 64706
rect 87950 64654 88002 64706
rect 97134 64654 97186 64706
rect 52446 64542 52498 64594
rect 56926 64542 56978 64594
rect 57486 64542 57538 64594
rect 57822 64542 57874 64594
rect 59390 64542 59442 64594
rect 60510 64542 60562 64594
rect 68574 64542 68626 64594
rect 69358 64542 69410 64594
rect 70478 64542 70530 64594
rect 71486 64542 71538 64594
rect 73278 64542 73330 64594
rect 75854 64542 75906 64594
rect 78206 64542 78258 64594
rect 78990 64542 79042 64594
rect 80894 64542 80946 64594
rect 84142 64542 84194 64594
rect 85374 64542 85426 64594
rect 86046 64542 86098 64594
rect 86270 64542 86322 64594
rect 86606 64542 86658 64594
rect 96350 64542 96402 64594
rect 52334 64430 52386 64482
rect 53566 64430 53618 64482
rect 55022 64430 55074 64482
rect 56366 64430 56418 64482
rect 56478 64430 56530 64482
rect 56702 64430 56754 64482
rect 57710 64430 57762 64482
rect 58494 64430 58546 64482
rect 58942 64430 58994 64482
rect 60286 64430 60338 64482
rect 74174 64430 74226 64482
rect 77198 64430 77250 64482
rect 77870 64430 77922 64482
rect 79326 64430 79378 64482
rect 80222 64430 80274 64482
rect 81118 64430 81170 64482
rect 82350 64430 82402 64482
rect 82910 64430 82962 64482
rect 83918 64430 83970 64482
rect 85150 64430 85202 64482
rect 86382 64430 86434 64482
rect 91198 64430 91250 64482
rect 93662 64430 93714 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 81278 64262 81330 64314
rect 81382 64262 81434 64314
rect 81486 64262 81538 64314
rect 58494 64094 58546 64146
rect 61630 64094 61682 64146
rect 66222 64094 66274 64146
rect 70926 64094 70978 64146
rect 72158 64094 72210 64146
rect 72718 64094 72770 64146
rect 74398 64094 74450 64146
rect 77646 64094 77698 64146
rect 78206 64094 78258 64146
rect 79326 64094 79378 64146
rect 79886 64094 79938 64146
rect 81902 64094 81954 64146
rect 82014 64094 82066 64146
rect 82910 64094 82962 64146
rect 83022 64094 83074 64146
rect 83134 64094 83186 64146
rect 85038 64094 85090 64146
rect 87054 64094 87106 64146
rect 87502 64094 87554 64146
rect 88398 64094 88450 64146
rect 90302 64094 90354 64146
rect 93438 64094 93490 64146
rect 94558 64094 94610 64146
rect 50318 63982 50370 64034
rect 54462 63982 54514 64034
rect 57486 63982 57538 64034
rect 66670 63982 66722 64034
rect 67678 63982 67730 64034
rect 70590 63982 70642 64034
rect 72382 63982 72434 64034
rect 73950 63982 74002 64034
rect 75966 63982 76018 64034
rect 77758 63982 77810 64034
rect 78430 63982 78482 64034
rect 80222 63982 80274 64034
rect 84814 63982 84866 64034
rect 96126 63982 96178 64034
rect 49534 63870 49586 63922
rect 52894 63870 52946 63922
rect 53902 63870 53954 63922
rect 54238 63870 54290 63922
rect 55134 63870 55186 63922
rect 55694 63870 55746 63922
rect 56590 63870 56642 63922
rect 57934 63870 57986 63922
rect 58270 63870 58322 63922
rect 59166 63870 59218 63922
rect 59726 63870 59778 63922
rect 60510 63870 60562 63922
rect 61182 63870 61234 63922
rect 67006 63870 67058 63922
rect 67454 63870 67506 63922
rect 68350 63870 68402 63922
rect 68798 63870 68850 63922
rect 69694 63870 69746 63922
rect 71374 63870 71426 63922
rect 71934 63870 71986 63922
rect 72606 63870 72658 63922
rect 75070 63870 75122 63922
rect 77086 63870 77138 63922
rect 77982 63870 78034 63922
rect 78990 63870 79042 63922
rect 81566 63870 81618 63922
rect 81790 63870 81842 63922
rect 82126 63870 82178 63922
rect 83246 63870 83298 63922
rect 83470 63870 83522 63922
rect 83918 63870 83970 63922
rect 85150 63870 85202 63922
rect 86046 63870 86098 63922
rect 86270 63870 86322 63922
rect 86606 63870 86658 63922
rect 89294 63870 89346 63922
rect 89630 63870 89682 63922
rect 90078 63870 90130 63922
rect 90750 63870 90802 63922
rect 91310 63870 91362 63922
rect 92318 63870 92370 63922
rect 92990 63870 93042 63922
rect 94334 63870 94386 63922
rect 96014 63870 96066 63922
rect 52446 63758 52498 63810
rect 53454 63758 53506 63810
rect 84366 63758 84418 63810
rect 86494 63758 86546 63810
rect 87950 63758 88002 63810
rect 95230 63646 95282 63698
rect 95566 63646 95618 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 96638 63478 96690 63530
rect 96742 63478 96794 63530
rect 96846 63478 96898 63530
rect 72046 63310 72098 63362
rect 50094 63198 50146 63250
rect 52222 63198 52274 63250
rect 52670 63198 52722 63250
rect 57486 63198 57538 63250
rect 58270 63198 58322 63250
rect 59502 63198 59554 63250
rect 66222 63198 66274 63250
rect 68126 63198 68178 63250
rect 77310 63198 77362 63250
rect 79326 63198 79378 63250
rect 86158 63198 86210 63250
rect 92206 63198 92258 63250
rect 96126 63198 96178 63250
rect 49422 63086 49474 63138
rect 54126 63086 54178 63138
rect 54462 63086 54514 63138
rect 55358 63086 55410 63138
rect 55694 63086 55746 63138
rect 56702 63086 56754 63138
rect 58158 63086 58210 63138
rect 58382 63086 58434 63138
rect 59390 63086 59442 63138
rect 59614 63086 59666 63138
rect 62414 63086 62466 63138
rect 67902 63086 67954 63138
rect 68238 63086 68290 63138
rect 68462 63086 68514 63138
rect 70142 63086 70194 63138
rect 71486 63086 71538 63138
rect 71934 63086 71986 63138
rect 72158 63086 72210 63138
rect 72718 63086 72770 63138
rect 76414 63086 76466 63138
rect 77758 63086 77810 63138
rect 78542 63086 78594 63138
rect 79662 63086 79714 63138
rect 80110 63086 80162 63138
rect 81006 63086 81058 63138
rect 81566 63086 81618 63138
rect 82350 63086 82402 63138
rect 83022 63086 83074 63138
rect 84254 63086 84306 63138
rect 86270 63086 86322 63138
rect 86494 63086 86546 63138
rect 88398 63086 88450 63138
rect 88846 63086 88898 63138
rect 89518 63086 89570 63138
rect 90078 63086 90130 63138
rect 91198 63086 91250 63138
rect 1822 62974 1874 63026
rect 53678 62974 53730 63026
rect 54686 62974 54738 63026
rect 58830 62974 58882 63026
rect 60062 62974 60114 63026
rect 61966 62974 62018 63026
rect 62302 62974 62354 63026
rect 67454 62974 67506 63026
rect 69246 62974 69298 63026
rect 73838 62974 73890 63026
rect 75854 62974 75906 63026
rect 78766 62974 78818 63026
rect 83582 62974 83634 63026
rect 83806 62974 83858 63026
rect 85822 62974 85874 63026
rect 86046 62974 86098 63026
rect 88062 62974 88114 63026
rect 94334 62974 94386 63026
rect 95006 62974 95058 63026
rect 95118 62974 95170 63026
rect 2158 62862 2210 62914
rect 58606 62862 58658 62914
rect 59838 62862 59890 62914
rect 62190 62862 62242 62914
rect 62974 62862 63026 62914
rect 63422 62862 63474 62914
rect 65886 62862 65938 62914
rect 67118 62862 67170 62914
rect 69806 62862 69858 62914
rect 70702 62862 70754 62914
rect 71710 62862 71762 62914
rect 76414 62862 76466 62914
rect 80334 62862 80386 62914
rect 83918 62862 83970 62914
rect 85150 62862 85202 62914
rect 86942 62862 86994 62914
rect 87390 62862 87442 62914
rect 89070 62862 89122 62914
rect 91758 62862 91810 62914
rect 93662 62862 93714 62914
rect 93998 62862 94050 62914
rect 94222 62862 94274 62914
rect 94782 62862 94834 62914
rect 95678 62862 95730 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 81278 62694 81330 62746
rect 81382 62694 81434 62746
rect 81486 62694 81538 62746
rect 56702 62526 56754 62578
rect 57598 62526 57650 62578
rect 59278 62526 59330 62578
rect 59502 62526 59554 62578
rect 60286 62526 60338 62578
rect 61966 62526 62018 62578
rect 63310 62526 63362 62578
rect 63982 62526 64034 62578
rect 75406 62526 75458 62578
rect 78430 62526 78482 62578
rect 81566 62526 81618 62578
rect 82462 62526 82514 62578
rect 84366 62526 84418 62578
rect 86270 62526 86322 62578
rect 86606 62526 86658 62578
rect 87614 62526 87666 62578
rect 90302 62526 90354 62578
rect 1822 62414 1874 62466
rect 48750 62414 48802 62466
rect 52670 62414 52722 62466
rect 57822 62414 57874 62466
rect 62190 62414 62242 62466
rect 62414 62414 62466 62466
rect 62974 62414 63026 62466
rect 63198 62414 63250 62466
rect 74846 62414 74898 62466
rect 77534 62414 77586 62466
rect 79438 62414 79490 62466
rect 79774 62414 79826 62466
rect 81342 62414 81394 62466
rect 81902 62414 81954 62466
rect 82798 62414 82850 62466
rect 84590 62414 84642 62466
rect 85150 62414 85202 62466
rect 87278 62414 87330 62466
rect 87502 62414 87554 62466
rect 87838 62414 87890 62466
rect 89294 62414 89346 62466
rect 90750 62414 90802 62466
rect 48414 62302 48466 62354
rect 55358 62302 55410 62354
rect 55806 62302 55858 62354
rect 57374 62302 57426 62354
rect 57934 62302 57986 62354
rect 58606 62302 58658 62354
rect 59166 62302 59218 62354
rect 61854 62302 61906 62354
rect 63534 62302 63586 62354
rect 66334 62302 66386 62354
rect 69918 62302 69970 62354
rect 70142 62302 70194 62354
rect 71038 62302 71090 62354
rect 72046 62302 72098 62354
rect 72494 62302 72546 62354
rect 75406 62302 75458 62354
rect 75742 62302 75794 62354
rect 78094 62302 78146 62354
rect 81678 62302 81730 62354
rect 83246 62302 83298 62354
rect 83694 62302 83746 62354
rect 84702 62302 84754 62354
rect 86046 62302 86098 62354
rect 86382 62302 86434 62354
rect 86494 62302 86546 62354
rect 89630 62302 89682 62354
rect 90190 62302 90242 62354
rect 91534 62302 91586 62354
rect 92318 62302 92370 62354
rect 93662 62302 93714 62354
rect 47854 62190 47906 62242
rect 59950 62190 60002 62242
rect 65774 62190 65826 62242
rect 67118 62190 67170 62242
rect 69246 62190 69298 62242
rect 71486 62190 71538 62242
rect 78878 62190 78930 62242
rect 80222 62190 80274 62242
rect 88286 62190 88338 62242
rect 93102 62190 93154 62242
rect 94334 62190 94386 62242
rect 96462 62190 96514 62242
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 96638 61910 96690 61962
rect 96742 61910 96794 61962
rect 96846 61910 96898 61962
rect 55134 61742 55186 61794
rect 70590 61742 70642 61794
rect 74174 61742 74226 61794
rect 82686 61742 82738 61794
rect 83134 61742 83186 61794
rect 48862 61630 48914 61682
rect 58606 61630 58658 61682
rect 65998 61630 66050 61682
rect 67902 61630 67954 61682
rect 68462 61630 68514 61682
rect 69246 61630 69298 61682
rect 71598 61630 71650 61682
rect 72494 61630 72546 61682
rect 74286 61630 74338 61682
rect 80446 61630 80498 61682
rect 82238 61630 82290 61682
rect 82686 61630 82738 61682
rect 83806 61630 83858 61682
rect 85710 61630 85762 61682
rect 86270 61630 86322 61682
rect 87614 61630 87666 61682
rect 88846 61630 88898 61682
rect 89182 61630 89234 61682
rect 93214 61630 93266 61682
rect 96798 61630 96850 61682
rect 49758 61518 49810 61570
rect 50430 61518 50482 61570
rect 58942 61518 58994 61570
rect 62302 61518 62354 61570
rect 62750 61518 62802 61570
rect 64094 61518 64146 61570
rect 64878 61518 64930 61570
rect 66558 61518 66610 61570
rect 67454 61518 67506 61570
rect 68126 61518 68178 61570
rect 70254 61518 70306 61570
rect 71150 61518 71202 61570
rect 72270 61518 72322 61570
rect 73950 61518 74002 61570
rect 74398 61518 74450 61570
rect 75182 61518 75234 61570
rect 75406 61518 75458 61570
rect 75630 61518 75682 61570
rect 75854 61518 75906 61570
rect 77310 61518 77362 61570
rect 78542 61518 78594 61570
rect 78990 61518 79042 61570
rect 79886 61518 79938 61570
rect 80670 61518 80722 61570
rect 80782 61518 80834 61570
rect 81678 61518 81730 61570
rect 83470 61518 83522 61570
rect 83694 61518 83746 61570
rect 85262 61518 85314 61570
rect 85486 61518 85538 61570
rect 85934 61518 85986 61570
rect 89630 61518 89682 61570
rect 93886 61518 93938 61570
rect 50318 61406 50370 61458
rect 55022 61406 55074 61458
rect 55694 61406 55746 61458
rect 59166 61406 59218 61458
rect 59278 61406 59330 61458
rect 60174 61406 60226 61458
rect 61854 61406 61906 61458
rect 62862 61406 62914 61458
rect 63310 61406 63362 61458
rect 67678 61406 67730 61458
rect 70030 61406 70082 61458
rect 70478 61406 70530 61458
rect 72830 61406 72882 61458
rect 79550 61406 79602 61458
rect 80334 61406 80386 61458
rect 81454 61406 81506 61458
rect 83918 61406 83970 61458
rect 94670 61406 94722 61458
rect 49422 61294 49474 61346
rect 51102 61294 51154 61346
rect 53342 61294 53394 61346
rect 55134 61294 55186 61346
rect 56142 61294 56194 61346
rect 59726 61294 59778 61346
rect 65550 61294 65602 61346
rect 66894 61294 66946 61346
rect 75966 61294 76018 61346
rect 76302 61294 76354 61346
rect 77870 61294 77922 61346
rect 79662 61294 79714 61346
rect 84366 61294 84418 61346
rect 86718 61294 86770 61346
rect 87166 61294 87218 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 81278 61126 81330 61178
rect 81382 61126 81434 61178
rect 81486 61126 81538 61178
rect 56254 60958 56306 61010
rect 62414 60958 62466 61010
rect 66670 60958 66722 61010
rect 69246 60958 69298 61010
rect 85822 60958 85874 61010
rect 88510 60958 88562 61010
rect 90638 60958 90690 61010
rect 48414 60846 48466 60898
rect 48750 60846 48802 60898
rect 50878 60846 50930 60898
rect 55470 60846 55522 60898
rect 65326 60846 65378 60898
rect 67230 60846 67282 60898
rect 68238 60846 68290 60898
rect 68574 60846 68626 60898
rect 70142 60846 70194 60898
rect 70478 60846 70530 60898
rect 71038 60846 71090 60898
rect 71374 60846 71426 60898
rect 72606 60846 72658 60898
rect 79326 60846 79378 60898
rect 79662 60846 79714 60898
rect 80558 60846 80610 60898
rect 82350 60846 82402 60898
rect 82798 60846 82850 60898
rect 84142 60846 84194 60898
rect 50094 60734 50146 60786
rect 50766 60734 50818 60786
rect 55246 60734 55298 60786
rect 55582 60734 55634 60786
rect 56142 60734 56194 60786
rect 56478 60734 56530 60786
rect 61854 60734 61906 60786
rect 62190 60734 62242 60786
rect 63086 60734 63138 60786
rect 63646 60734 63698 60786
rect 64542 60734 64594 60786
rect 67566 60734 67618 60786
rect 69358 60734 69410 60786
rect 72158 60734 72210 60786
rect 78766 60734 78818 60786
rect 80222 60734 80274 60786
rect 81342 60734 81394 60786
rect 83246 60734 83298 60786
rect 84254 60734 84306 60786
rect 85150 60734 85202 60786
rect 85598 60734 85650 60786
rect 86382 60734 86434 60786
rect 87054 60734 87106 60786
rect 87950 60734 88002 60786
rect 89742 60734 89794 60786
rect 95790 60734 95842 60786
rect 51438 60622 51490 60674
rect 51886 60622 51938 60674
rect 57374 60622 57426 60674
rect 57822 60622 57874 60674
rect 61406 60622 61458 60674
rect 65886 60622 65938 60674
rect 66222 60622 66274 60674
rect 76750 60622 76802 60674
rect 81902 60622 81954 60674
rect 84814 60622 84866 60674
rect 89294 60622 89346 60674
rect 93550 60622 93602 60674
rect 49758 60510 49810 60562
rect 65886 60510 65938 60562
rect 66558 60510 66610 60562
rect 69246 60510 69298 60562
rect 81454 60510 81506 60562
rect 84142 60510 84194 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 96638 60342 96690 60394
rect 96742 60342 96794 60394
rect 96846 60342 96898 60394
rect 57262 60174 57314 60226
rect 66110 60174 66162 60226
rect 66782 60174 66834 60226
rect 72718 60174 72770 60226
rect 72942 60174 72994 60226
rect 74958 60174 75010 60226
rect 49086 60062 49138 60114
rect 51214 60062 51266 60114
rect 56590 60062 56642 60114
rect 67230 60062 67282 60114
rect 68462 60062 68514 60114
rect 71486 60062 71538 60114
rect 75854 60062 75906 60114
rect 83134 60062 83186 60114
rect 83582 60062 83634 60114
rect 84030 60062 84082 60114
rect 89070 60062 89122 60114
rect 96462 60062 96514 60114
rect 48414 59950 48466 60002
rect 51774 59950 51826 60002
rect 52782 59950 52834 60002
rect 53678 59950 53730 60002
rect 62862 59950 62914 60002
rect 63646 59950 63698 60002
rect 64430 59950 64482 60002
rect 65102 59950 65154 60002
rect 65550 59950 65602 60002
rect 67678 59950 67730 60002
rect 68014 59950 68066 60002
rect 69470 59950 69522 60002
rect 71934 59950 71986 60002
rect 72494 59950 72546 60002
rect 73950 59950 74002 60002
rect 74510 59950 74562 60002
rect 75294 59950 75346 60002
rect 79774 59950 79826 60002
rect 80222 59950 80274 60002
rect 80894 59950 80946 60002
rect 81678 59950 81730 60002
rect 82462 59950 82514 60002
rect 85598 59950 85650 60002
rect 86046 59950 86098 60002
rect 87502 59950 87554 60002
rect 88398 59950 88450 60002
rect 92206 59950 92258 60002
rect 92542 59950 92594 60002
rect 93550 59950 93602 60002
rect 94334 59950 94386 60002
rect 97694 59950 97746 60002
rect 54462 59838 54514 59890
rect 57262 59838 57314 59890
rect 57374 59838 57426 59890
rect 58382 59838 58434 59890
rect 58494 59838 58546 59890
rect 64878 59838 64930 59890
rect 65886 59838 65938 59890
rect 66782 59838 66834 59890
rect 69806 59838 69858 59890
rect 70478 59838 70530 59890
rect 70814 59838 70866 59890
rect 73054 59838 73106 59890
rect 74062 59838 74114 59890
rect 76414 59838 76466 59890
rect 77646 59838 77698 59890
rect 78206 59838 78258 59890
rect 78542 59838 78594 59890
rect 79438 59838 79490 59890
rect 80446 59838 80498 59890
rect 84478 59838 84530 59890
rect 85262 59838 85314 59890
rect 86270 59838 86322 59890
rect 86718 59838 86770 59890
rect 97022 59838 97074 59890
rect 97134 59838 97186 59890
rect 97358 59838 97410 59890
rect 98030 59838 98082 59890
rect 58158 59726 58210 59778
rect 58942 59726 58994 59778
rect 61742 59726 61794 59778
rect 62190 59726 62242 59778
rect 66334 59726 66386 59778
rect 67902 59726 67954 59778
rect 77310 59726 77362 59778
rect 89406 59726 89458 59778
rect 89854 59726 89906 59778
rect 92318 59726 92370 59778
rect 97918 59726 97970 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 81278 59558 81330 59610
rect 81382 59558 81434 59610
rect 81486 59558 81538 59610
rect 48750 59390 48802 59442
rect 58158 59390 58210 59442
rect 63870 59390 63922 59442
rect 67902 59390 67954 59442
rect 70590 59390 70642 59442
rect 71150 59390 71202 59442
rect 75518 59390 75570 59442
rect 80334 59390 80386 59442
rect 81230 59390 81282 59442
rect 82126 59390 82178 59442
rect 83134 59390 83186 59442
rect 83470 59390 83522 59442
rect 84366 59390 84418 59442
rect 94222 59390 94274 59442
rect 97134 59390 97186 59442
rect 47854 59278 47906 59330
rect 50318 59278 50370 59330
rect 54574 59278 54626 59330
rect 57598 59278 57650 59330
rect 58382 59278 58434 59330
rect 58494 59278 58546 59330
rect 63086 59278 63138 59330
rect 69358 59278 69410 59330
rect 74398 59278 74450 59330
rect 76974 59278 77026 59330
rect 78094 59278 78146 59330
rect 78990 59278 79042 59330
rect 89630 59278 89682 59330
rect 94446 59278 94498 59330
rect 94558 59278 94610 59330
rect 95566 59278 95618 59330
rect 95790 59278 95842 59330
rect 46958 59166 47010 59218
rect 47630 59166 47682 59218
rect 48526 59166 48578 59218
rect 49534 59166 49586 59218
rect 53790 59166 53842 59218
rect 57710 59166 57762 59218
rect 59614 59166 59666 59218
rect 62862 59166 62914 59218
rect 63198 59166 63250 59218
rect 63646 59166 63698 59218
rect 63982 59166 64034 59218
rect 65886 59166 65938 59218
rect 66894 59166 66946 59218
rect 67342 59166 67394 59218
rect 68126 59166 68178 59218
rect 68574 59166 68626 59218
rect 70366 59166 70418 59218
rect 71374 59166 71426 59218
rect 72046 59166 72098 59218
rect 72606 59166 72658 59218
rect 75518 59166 75570 59218
rect 75854 59166 75906 59218
rect 78430 59166 78482 59218
rect 79326 59166 79378 59218
rect 89518 59166 89570 59218
rect 89854 59166 89906 59218
rect 95902 59166 95954 59218
rect 52446 59054 52498 59106
rect 53006 59054 53058 59106
rect 56702 59054 56754 59106
rect 58942 59054 58994 59106
rect 60286 59054 60338 59106
rect 62414 59054 62466 59106
rect 64542 59054 64594 59106
rect 68910 59054 68962 59106
rect 78206 59054 78258 59106
rect 79774 59054 79826 59106
rect 81678 59054 81730 59106
rect 82574 59054 82626 59106
rect 83918 59054 83970 59106
rect 84814 59054 84866 59106
rect 85262 59054 85314 59106
rect 85710 59054 85762 59106
rect 91758 59054 91810 59106
rect 96350 59054 96402 59106
rect 57598 58942 57650 58994
rect 82462 58942 82514 58994
rect 83918 58942 83970 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 96638 58774 96690 58826
rect 96742 58774 96794 58826
rect 96846 58774 96898 58826
rect 51102 58606 51154 58658
rect 51662 58606 51714 58658
rect 64990 58606 65042 58658
rect 69134 58606 69186 58658
rect 69806 58606 69858 58658
rect 83470 58606 83522 58658
rect 84478 58606 84530 58658
rect 47966 58494 48018 58546
rect 51102 58494 51154 58546
rect 51998 58494 52050 58546
rect 58046 58494 58098 58546
rect 61406 58494 61458 58546
rect 63534 58494 63586 58546
rect 69358 58494 69410 58546
rect 70254 58494 70306 58546
rect 72270 58494 72322 58546
rect 78878 58494 78930 58546
rect 80222 58494 80274 58546
rect 81118 58494 81170 58546
rect 83134 58494 83186 58546
rect 83582 58494 83634 58546
rect 84142 58494 84194 58546
rect 84478 58494 84530 58546
rect 85150 58494 85202 58546
rect 88510 58494 88562 58546
rect 90638 58494 90690 58546
rect 48526 58382 48578 58434
rect 49422 58382 49474 58434
rect 49758 58382 49810 58434
rect 50542 58382 50594 58434
rect 54350 58382 54402 58434
rect 55246 58382 55298 58434
rect 58494 58382 58546 58434
rect 59838 58382 59890 58434
rect 60286 58382 60338 58434
rect 64206 58382 64258 58434
rect 65102 58382 65154 58434
rect 68238 58382 68290 58434
rect 68574 58382 68626 58434
rect 72158 58382 72210 58434
rect 73502 58382 73554 58434
rect 74062 58382 74114 58434
rect 74622 58382 74674 58434
rect 75630 58382 75682 58434
rect 76078 58382 76130 58434
rect 79774 58382 79826 58434
rect 91422 58382 91474 58434
rect 95678 58382 95730 58434
rect 50430 58270 50482 58322
rect 54462 58270 54514 58322
rect 54686 58270 54738 58322
rect 55918 58270 55970 58322
rect 60622 58270 60674 58322
rect 65550 58270 65602 58322
rect 65774 58270 65826 58322
rect 65886 58270 65938 58322
rect 70814 58270 70866 58322
rect 71150 58270 71202 58322
rect 71822 58270 71874 58322
rect 73278 58270 73330 58322
rect 73614 58270 73666 58322
rect 75406 58270 75458 58322
rect 77310 58270 77362 58322
rect 77646 58270 77698 58322
rect 78206 58270 78258 58322
rect 78318 58270 78370 58322
rect 81566 58270 81618 58322
rect 87726 58270 87778 58322
rect 87838 58270 87890 58322
rect 94894 58270 94946 58322
rect 96462 58270 96514 58322
rect 48750 58158 48802 58210
rect 51662 58158 51714 58210
rect 52670 58158 52722 58210
rect 53454 58158 53506 58210
rect 60510 58158 60562 58210
rect 64990 58158 65042 58210
rect 66446 58158 66498 58210
rect 66894 58158 66946 58210
rect 69806 58158 69858 58210
rect 72830 58158 72882 58210
rect 75294 58158 75346 58210
rect 75854 58158 75906 58210
rect 76526 58158 76578 58210
rect 78542 58158 78594 58210
rect 79326 58158 79378 58210
rect 80670 58158 80722 58210
rect 82126 58158 82178 58210
rect 86830 58158 86882 58210
rect 87278 58158 87330 58210
rect 88062 58158 88114 58210
rect 91982 58158 92034 58210
rect 92430 58158 92482 58210
rect 93214 58158 93266 58210
rect 94558 58158 94610 58210
rect 94782 58158 94834 58210
rect 95342 58158 95394 58210
rect 95566 58158 95618 58210
rect 96126 58158 96178 58210
rect 96350 58158 96402 58210
rect 96910 58158 96962 58210
rect 97358 58158 97410 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 81278 57990 81330 58042
rect 81382 57990 81434 58042
rect 81486 57990 81538 58042
rect 51438 57822 51490 57874
rect 65326 57822 65378 57874
rect 65550 57822 65602 57874
rect 66110 57822 66162 57874
rect 69582 57822 69634 57874
rect 70030 57822 70082 57874
rect 70366 57822 70418 57874
rect 73502 57822 73554 57874
rect 76190 57822 76242 57874
rect 77422 57822 77474 57874
rect 78878 57822 78930 57874
rect 82014 57822 82066 57874
rect 97582 57822 97634 57874
rect 50654 57710 50706 57762
rect 53118 57710 53170 57762
rect 57598 57710 57650 57762
rect 57710 57710 57762 57762
rect 60958 57710 61010 57762
rect 65662 57710 65714 57762
rect 73614 57710 73666 57762
rect 74846 57710 74898 57762
rect 75854 57710 75906 57762
rect 76862 57710 76914 57762
rect 76974 57710 77026 57762
rect 78542 57710 78594 57762
rect 79438 57710 79490 57762
rect 79550 57710 79602 57762
rect 80334 57710 80386 57762
rect 80446 57710 80498 57762
rect 80670 57710 80722 57762
rect 81342 57710 81394 57762
rect 81454 57710 81506 57762
rect 84702 57710 84754 57762
rect 88286 57710 88338 57762
rect 88398 57710 88450 57762
rect 92766 57710 92818 57762
rect 92878 57710 92930 57762
rect 94334 57710 94386 57762
rect 97246 57710 97298 57762
rect 97358 57710 97410 57762
rect 50766 57598 50818 57650
rect 51774 57598 51826 57650
rect 53006 57598 53058 57650
rect 53342 57598 53394 57650
rect 53790 57598 53842 57650
rect 60398 57598 60450 57650
rect 67006 57598 67058 57650
rect 67566 57598 67618 57650
rect 71598 57598 71650 57650
rect 71822 57598 71874 57650
rect 74286 57598 74338 57650
rect 74734 57598 74786 57650
rect 75070 57598 75122 57650
rect 75742 57598 75794 57650
rect 82910 57598 82962 57650
rect 84030 57598 84082 57650
rect 84478 57598 84530 57650
rect 85262 57598 85314 57650
rect 85934 57598 85986 57650
rect 86830 57598 86882 57650
rect 88622 57598 88674 57650
rect 91422 57598 91474 57650
rect 92206 57598 92258 57650
rect 93102 57598 93154 57650
rect 93662 57598 93714 57650
rect 52222 57486 52274 57538
rect 54574 57486 54626 57538
rect 56702 57486 56754 57538
rect 64766 57486 64818 57538
rect 68014 57486 68066 57538
rect 68798 57486 68850 57538
rect 70814 57486 70866 57538
rect 72606 57486 72658 57538
rect 77870 57486 77922 57538
rect 82574 57486 82626 57538
rect 83694 57486 83746 57538
rect 87502 57486 87554 57538
rect 89294 57486 89346 57538
rect 96462 57486 96514 57538
rect 97918 57486 97970 57538
rect 49646 57374 49698 57426
rect 49982 57374 50034 57426
rect 57598 57374 57650 57426
rect 72158 57374 72210 57426
rect 73502 57374 73554 57426
rect 74062 57374 74114 57426
rect 79550 57374 79602 57426
rect 81454 57374 81506 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 96638 57206 96690 57258
rect 96742 57206 96794 57258
rect 96846 57206 96898 57258
rect 57374 57038 57426 57090
rect 88622 57038 88674 57090
rect 49086 56926 49138 56978
rect 51214 56926 51266 56978
rect 54350 56926 54402 56978
rect 56478 56926 56530 56978
rect 62190 56926 62242 56978
rect 64318 56926 64370 56978
rect 70142 56926 70194 56978
rect 70590 56926 70642 56978
rect 72718 56926 72770 56978
rect 73054 56926 73106 56978
rect 73614 56926 73666 56978
rect 76414 56926 76466 56978
rect 78990 56926 79042 56978
rect 81118 56926 81170 56978
rect 87390 56926 87442 56978
rect 87950 56926 88002 56978
rect 92206 56926 92258 56978
rect 95006 56926 95058 56978
rect 97134 56926 97186 56978
rect 48414 56814 48466 56866
rect 53566 56814 53618 56866
rect 57486 56814 57538 56866
rect 57934 56814 57986 56866
rect 61518 56814 61570 56866
rect 68126 56814 68178 56866
rect 68574 56814 68626 56866
rect 69694 56814 69746 56866
rect 71822 56814 71874 56866
rect 73838 56814 73890 56866
rect 74174 56814 74226 56866
rect 78206 56814 78258 56866
rect 81566 56814 81618 56866
rect 83246 56814 83298 56866
rect 84030 56814 84082 56866
rect 88510 56814 88562 56866
rect 89406 56814 89458 56866
rect 93438 56814 93490 56866
rect 94334 56814 94386 56866
rect 57374 56702 57426 56754
rect 58270 56702 58322 56754
rect 74958 56702 75010 56754
rect 75294 56702 75346 56754
rect 75966 56702 76018 56754
rect 81790 56702 81842 56754
rect 81902 56702 81954 56754
rect 83470 56702 83522 56754
rect 88622 56702 88674 56754
rect 90078 56702 90130 56754
rect 51662 56590 51714 56642
rect 52670 56590 52722 56642
rect 58158 56590 58210 56642
rect 58718 56590 58770 56642
rect 59166 56590 59218 56642
rect 64766 56590 64818 56642
rect 65214 56590 65266 56642
rect 69358 56590 69410 56642
rect 71150 56590 71202 56642
rect 71598 56590 71650 56642
rect 75854 56590 75906 56642
rect 77198 56590 77250 56642
rect 77646 56590 77698 56642
rect 82574 56590 82626 56642
rect 84366 56590 84418 56642
rect 85150 56590 85202 56642
rect 93102 56590 93154 56642
rect 93326 56590 93378 56642
rect 97582 56590 97634 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 81278 56422 81330 56474
rect 81382 56422 81434 56474
rect 81486 56422 81538 56474
rect 50654 56254 50706 56306
rect 57374 56254 57426 56306
rect 68014 56254 68066 56306
rect 68238 56254 68290 56306
rect 70926 56254 70978 56306
rect 71486 56254 71538 56306
rect 71934 56254 71986 56306
rect 72494 56254 72546 56306
rect 73726 56254 73778 56306
rect 73950 56254 74002 56306
rect 75406 56254 75458 56306
rect 77310 56254 77362 56306
rect 77870 56254 77922 56306
rect 79438 56254 79490 56306
rect 80334 56254 80386 56306
rect 88622 56254 88674 56306
rect 90526 56254 90578 56306
rect 51438 56142 51490 56194
rect 57598 56142 57650 56194
rect 57710 56142 57762 56194
rect 60846 56142 60898 56194
rect 60958 56142 61010 56194
rect 65550 56142 65602 56194
rect 67454 56142 67506 56194
rect 67566 56142 67618 56194
rect 72382 56142 72434 56194
rect 73502 56142 73554 56194
rect 74510 56142 74562 56194
rect 74846 56142 74898 56194
rect 76302 56142 76354 56194
rect 76638 56142 76690 56194
rect 77422 56142 77474 56194
rect 78878 56142 78930 56194
rect 79998 56142 80050 56194
rect 88286 56142 88338 56194
rect 88398 56142 88450 56194
rect 89630 56142 89682 56194
rect 89742 56142 89794 56194
rect 90302 56142 90354 56194
rect 56478 56030 56530 56082
rect 61630 56030 61682 56082
rect 65326 56030 65378 56082
rect 65662 56030 65714 56082
rect 66110 56030 66162 56082
rect 68350 56030 68402 56082
rect 68910 56030 68962 56082
rect 75742 56030 75794 56082
rect 77086 56030 77138 56082
rect 78766 56030 78818 56082
rect 82798 56030 82850 56082
rect 87502 56030 87554 56082
rect 90638 56030 90690 56082
rect 92318 56030 92370 56082
rect 58158 55918 58210 55970
rect 62414 55918 62466 55970
rect 64542 55918 64594 55970
rect 84030 55918 84082 55970
rect 96238 55918 96290 55970
rect 97246 55918 97298 55970
rect 60958 55806 61010 55858
rect 67454 55806 67506 55858
rect 72494 55806 72546 55858
rect 74062 55806 74114 55858
rect 78878 55806 78930 55858
rect 89742 55806 89794 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 96638 55638 96690 55690
rect 96742 55638 96794 55690
rect 96846 55638 96898 55690
rect 78990 55470 79042 55522
rect 51214 55358 51266 55410
rect 54462 55358 54514 55410
rect 56590 55358 56642 55410
rect 80558 55358 80610 55410
rect 82686 55358 82738 55410
rect 88174 55358 88226 55410
rect 89742 55358 89794 55410
rect 91870 55358 91922 55410
rect 92318 55358 92370 55410
rect 94334 55358 94386 55410
rect 96462 55358 96514 55410
rect 96910 55358 96962 55410
rect 48414 55246 48466 55298
rect 53790 55246 53842 55298
rect 60622 55246 60674 55298
rect 68574 55246 68626 55298
rect 70702 55246 70754 55298
rect 72046 55246 72098 55298
rect 72718 55246 72770 55298
rect 74958 55246 75010 55298
rect 77758 55246 77810 55298
rect 78318 55246 78370 55298
rect 79774 55246 79826 55298
rect 83358 55246 83410 55298
rect 84366 55246 84418 55298
rect 85262 55246 85314 55298
rect 89070 55246 89122 55298
rect 93550 55246 93602 55298
rect 49086 55134 49138 55186
rect 51774 55134 51826 55186
rect 52110 55134 52162 55186
rect 52558 55134 52610 55186
rect 61294 55134 61346 55186
rect 62414 55134 62466 55186
rect 63870 55134 63922 55186
rect 73390 55134 73442 55186
rect 76526 55134 76578 55186
rect 77198 55134 77250 55186
rect 78990 55134 79042 55186
rect 57038 55022 57090 55074
rect 62078 55022 62130 55074
rect 62302 55022 62354 55074
rect 68574 55022 68626 55074
rect 68798 55022 68850 55074
rect 70926 55022 70978 55074
rect 79102 55078 79154 55130
rect 83582 55134 83634 55186
rect 86046 55134 86098 55186
rect 71822 55022 71874 55074
rect 75518 55022 75570 55074
rect 84142 55022 84194 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 81278 54854 81330 54906
rect 81382 54854 81434 54906
rect 81486 54854 81538 54906
rect 48750 54686 48802 54738
rect 54350 54686 54402 54738
rect 55470 54686 55522 54738
rect 56702 54686 56754 54738
rect 59726 54686 59778 54738
rect 63982 54686 64034 54738
rect 72270 54686 72322 54738
rect 72606 54686 72658 54738
rect 74958 54686 75010 54738
rect 85598 54686 85650 54738
rect 86046 54686 86098 54738
rect 87502 54686 87554 54738
rect 88510 54686 88562 54738
rect 89294 54686 89346 54738
rect 90862 54686 90914 54738
rect 93102 54686 93154 54738
rect 93886 54686 93938 54738
rect 94670 54686 94722 54738
rect 48414 54574 48466 54626
rect 50878 54574 50930 54626
rect 52894 54574 52946 54626
rect 55694 54574 55746 54626
rect 56478 54574 56530 54626
rect 59950 54574 60002 54626
rect 61406 54574 61458 54626
rect 64206 54574 64258 54626
rect 64318 54574 64370 54626
rect 66446 54574 66498 54626
rect 69134 54574 69186 54626
rect 69470 54574 69522 54626
rect 69918 54574 69970 54626
rect 71150 54574 71202 54626
rect 76414 54574 76466 54626
rect 76750 54574 76802 54626
rect 78430 54574 78482 54626
rect 82574 54574 82626 54626
rect 85262 54574 85314 54626
rect 88286 54574 88338 54626
rect 89518 54574 89570 54626
rect 90302 54574 90354 54626
rect 91086 54574 91138 54626
rect 92766 54574 92818 54626
rect 92878 54574 92930 54626
rect 93550 54574 93602 54626
rect 93662 54574 93714 54626
rect 94446 54574 94498 54626
rect 50206 54462 50258 54514
rect 50990 54462 51042 54514
rect 52110 54462 52162 54514
rect 52782 54462 52834 54514
rect 55022 54462 55074 54514
rect 55806 54462 55858 54514
rect 56366 54462 56418 54514
rect 60062 54462 60114 54514
rect 60734 54462 60786 54514
rect 65662 54462 65714 54514
rect 73838 54462 73890 54514
rect 74062 54462 74114 54514
rect 77758 54462 77810 54514
rect 81790 54462 81842 54514
rect 86830 54462 86882 54514
rect 87390 54462 87442 54514
rect 88174 54462 88226 54514
rect 89630 54462 89682 54514
rect 90078 54462 90130 54514
rect 90414 54462 90466 54514
rect 91198 54462 91250 54514
rect 94334 54462 94386 54514
rect 53454 54350 53506 54402
rect 53902 54350 53954 54402
rect 57374 54350 57426 54402
rect 57822 54350 57874 54402
rect 59278 54350 59330 54402
rect 63534 54350 63586 54402
rect 68574 54350 68626 54402
rect 71710 54350 71762 54402
rect 73390 54350 73442 54402
rect 75406 54350 75458 54402
rect 80558 54350 80610 54402
rect 81342 54350 81394 54402
rect 84702 54350 84754 54402
rect 91646 54350 91698 54402
rect 92094 54350 92146 54402
rect 95006 54350 95058 54402
rect 98030 54350 98082 54402
rect 49870 54238 49922 54290
rect 51774 54238 51826 54290
rect 73614 54238 73666 54290
rect 74510 54238 74562 54290
rect 87502 54238 87554 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 96638 54070 96690 54122
rect 96742 54070 96794 54122
rect 96846 54070 96898 54122
rect 60062 53902 60114 53954
rect 60286 53902 60338 53954
rect 72606 53902 72658 53954
rect 73614 53902 73666 53954
rect 83806 53902 83858 53954
rect 84142 53902 84194 53954
rect 51662 53790 51714 53842
rect 64318 53790 64370 53842
rect 74734 53790 74786 53842
rect 75854 53790 75906 53842
rect 80222 53790 80274 53842
rect 87838 53790 87890 53842
rect 91646 53790 91698 53842
rect 93102 53790 93154 53842
rect 93662 53790 93714 53842
rect 94110 53790 94162 53842
rect 94782 53790 94834 53842
rect 47966 53678 48018 53730
rect 48862 53678 48914 53730
rect 52110 53678 52162 53730
rect 56366 53678 56418 53730
rect 56702 53678 56754 53730
rect 57486 53678 57538 53730
rect 61518 53678 61570 53730
rect 62190 53678 62242 53730
rect 64766 53678 64818 53730
rect 65326 53678 65378 53730
rect 67006 53678 67058 53730
rect 67454 53678 67506 53730
rect 67790 53678 67842 53730
rect 76302 53678 76354 53730
rect 77422 53678 77474 53730
rect 83246 53678 83298 53730
rect 87278 53678 87330 53730
rect 90750 53678 90802 53730
rect 91198 53678 91250 53730
rect 92318 53678 92370 53730
rect 97694 53678 97746 53730
rect 48190 53566 48242 53618
rect 49534 53566 49586 53618
rect 65550 53566 65602 53618
rect 65662 53566 65714 53618
rect 66110 53566 66162 53618
rect 68574 53566 68626 53618
rect 69582 53566 69634 53618
rect 70366 53566 70418 53618
rect 76414 53566 76466 53618
rect 76638 53566 76690 53618
rect 78094 53566 78146 53618
rect 83022 53566 83074 53618
rect 85150 53566 85202 53618
rect 86382 53566 86434 53618
rect 86942 53566 86994 53618
rect 89966 53566 90018 53618
rect 96910 53566 96962 53618
rect 52558 53454 52610 53506
rect 56478 53454 56530 53506
rect 57150 53454 57202 53506
rect 60286 53454 60338 53506
rect 67678 53454 67730 53506
rect 68238 53454 68290 53506
rect 68462 53454 68514 53506
rect 69246 53454 69298 53506
rect 69470 53454 69522 53506
rect 70030 53454 70082 53506
rect 70254 53454 70306 53506
rect 70814 53454 70866 53506
rect 71262 53454 71314 53506
rect 72494 53454 72546 53506
rect 73054 53454 73106 53506
rect 73502 53454 73554 53506
rect 80670 53454 80722 53506
rect 82350 53454 82402 53506
rect 87054 53454 87106 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 81278 53286 81330 53338
rect 81382 53286 81434 53338
rect 81486 53286 81538 53338
rect 52894 53118 52946 53170
rect 61630 53118 61682 53170
rect 61854 53118 61906 53170
rect 62862 53118 62914 53170
rect 63198 53118 63250 53170
rect 63422 53118 63474 53170
rect 65326 53118 65378 53170
rect 65774 53118 65826 53170
rect 70366 53118 70418 53170
rect 71150 53118 71202 53170
rect 72270 53118 72322 53170
rect 75294 53118 75346 53170
rect 75742 53118 75794 53170
rect 77646 53118 77698 53170
rect 78430 53118 78482 53170
rect 78654 53118 78706 53170
rect 79550 53118 79602 53170
rect 83022 53118 83074 53170
rect 89406 53118 89458 53170
rect 89630 53118 89682 53170
rect 90526 53118 90578 53170
rect 92206 53118 92258 53170
rect 95678 53118 95730 53170
rect 98030 53118 98082 53170
rect 62638 53006 62690 53058
rect 63534 53006 63586 53058
rect 64542 53006 64594 53058
rect 67342 53006 67394 53058
rect 70814 53006 70866 53058
rect 87390 53006 87442 53058
rect 89294 53006 89346 53058
rect 94670 53006 94722 53058
rect 95454 53006 95506 53058
rect 96238 53006 96290 53058
rect 49534 52894 49586 52946
rect 61966 52894 62018 52946
rect 62526 52894 62578 52946
rect 66558 52894 66610 52946
rect 73390 52894 73442 52946
rect 78318 52894 78370 52946
rect 79102 52894 79154 52946
rect 88174 52894 88226 52946
rect 90078 52894 90130 52946
rect 94558 52894 94610 52946
rect 95342 52894 95394 52946
rect 96126 52894 96178 52946
rect 96462 52894 96514 52946
rect 97582 52894 97634 52946
rect 50318 52782 50370 52834
rect 52446 52782 52498 52834
rect 61182 52782 61234 52834
rect 63982 52782 64034 52834
rect 69470 52782 69522 52834
rect 71710 52782 71762 52834
rect 73838 52782 73890 52834
rect 74398 52782 74450 52834
rect 85262 52782 85314 52834
rect 90862 52782 90914 52834
rect 92654 52782 92706 52834
rect 93214 52782 93266 52834
rect 93550 52782 93602 52834
rect 93998 52782 94050 52834
rect 97134 52782 97186 52834
rect 94670 52670 94722 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 96638 52502 96690 52554
rect 96742 52502 96794 52554
rect 96846 52502 96898 52554
rect 62190 52334 62242 52386
rect 62638 52334 62690 52386
rect 53342 52222 53394 52274
rect 62190 52222 62242 52274
rect 66334 52222 66386 52274
rect 69806 52222 69858 52274
rect 73502 52222 73554 52274
rect 73950 52222 74002 52274
rect 77646 52222 77698 52274
rect 78766 52222 78818 52274
rect 86046 52222 86098 52274
rect 94782 52222 94834 52274
rect 53790 52110 53842 52162
rect 54574 52110 54626 52162
rect 55022 52110 55074 52162
rect 55358 52110 55410 52162
rect 56254 52110 56306 52162
rect 56590 52110 56642 52162
rect 57598 52110 57650 52162
rect 58718 52110 58770 52162
rect 62638 52110 62690 52162
rect 67006 52110 67058 52162
rect 68126 52110 68178 52162
rect 70142 52110 70194 52162
rect 70702 52110 70754 52162
rect 71262 52110 71314 52162
rect 72046 52110 72098 52162
rect 72830 52110 72882 52162
rect 74734 52110 74786 52162
rect 75742 52110 75794 52162
rect 76302 52110 76354 52162
rect 85486 52110 85538 52162
rect 86382 52110 86434 52162
rect 86942 52110 86994 52162
rect 87502 52110 87554 52162
rect 88286 52110 88338 52162
rect 89182 52110 89234 52162
rect 91198 52110 91250 52162
rect 92430 52110 92482 52162
rect 94334 52110 94386 52162
rect 97694 52110 97746 52162
rect 49310 51998 49362 52050
rect 49646 51998 49698 52050
rect 55582 51998 55634 52050
rect 67118 51998 67170 52050
rect 67790 51998 67842 52050
rect 67902 51998 67954 52050
rect 68462 51998 68514 52050
rect 70814 51998 70866 52050
rect 87054 51998 87106 52050
rect 89854 51998 89906 52050
rect 93326 51998 93378 52050
rect 93438 51998 93490 52050
rect 93998 51998 94050 52050
rect 94110 51998 94162 52050
rect 96910 51998 96962 52050
rect 58270 51886 58322 51938
rect 67342 51886 67394 51938
rect 75070 51886 75122 51938
rect 77198 51886 77250 51938
rect 90190 51886 90242 51938
rect 91422 51886 91474 51938
rect 91870 51886 91922 51938
rect 93102 51886 93154 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 81278 51718 81330 51770
rect 81382 51718 81434 51770
rect 81486 51718 81538 51770
rect 53118 51550 53170 51602
rect 54350 51550 54402 51602
rect 57374 51550 57426 51602
rect 60174 51550 60226 51602
rect 61630 51550 61682 51602
rect 62078 51550 62130 51602
rect 63982 51550 64034 51602
rect 65326 51550 65378 51602
rect 74062 51550 74114 51602
rect 74510 51550 74562 51602
rect 75518 51550 75570 51602
rect 76862 51550 76914 51602
rect 77422 51550 77474 51602
rect 82462 51550 82514 51602
rect 89630 51550 89682 51602
rect 97134 51550 97186 51602
rect 97358 51550 97410 51602
rect 97918 51550 97970 51602
rect 59726 51438 59778 51490
rect 68014 51438 68066 51490
rect 73502 51438 73554 51490
rect 75854 51438 75906 51490
rect 78318 51438 78370 51490
rect 79102 51438 79154 51490
rect 79214 51438 79266 51490
rect 79438 51438 79490 51490
rect 79998 51438 80050 51490
rect 81230 51438 81282 51490
rect 81454 51438 81506 51490
rect 96238 51438 96290 51490
rect 97470 51438 97522 51490
rect 58046 51326 58098 51378
rect 59166 51326 59218 51378
rect 60286 51326 60338 51378
rect 60846 51326 60898 51378
rect 64094 51326 64146 51378
rect 67342 51326 67394 51378
rect 73278 51326 73330 51378
rect 73614 51326 73666 51378
rect 76750 51326 76802 51378
rect 77086 51326 77138 51378
rect 78206 51326 78258 51378
rect 79886 51326 79938 51378
rect 81566 51326 81618 51378
rect 91982 51326 92034 51378
rect 54798 51214 54850 51266
rect 55246 51214 55298 51266
rect 55694 51214 55746 51266
rect 56030 51214 56082 51266
rect 61182 51214 61234 51266
rect 62638 51214 62690 51266
rect 62974 51214 63026 51266
rect 64542 51214 64594 51266
rect 70142 51214 70194 51266
rect 70702 51214 70754 51266
rect 71038 51214 71090 51266
rect 71710 51214 71762 51266
rect 75070 51214 75122 51266
rect 80558 51214 80610 51266
rect 82014 51214 82066 51266
rect 85710 51214 85762 51266
rect 89966 51214 90018 51266
rect 90414 51214 90466 51266
rect 54238 51102 54290 51154
rect 55246 51102 55298 51154
rect 63982 51102 64034 51154
rect 78318 51102 78370 51154
rect 79998 51102 80050 51154
rect 89518 51102 89570 51154
rect 90414 51102 90466 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 96638 50934 96690 50986
rect 96742 50934 96794 50986
rect 96846 50934 96898 50986
rect 65998 50766 66050 50818
rect 66558 50766 66610 50818
rect 93326 50766 93378 50818
rect 58382 50654 58434 50706
rect 58942 50654 58994 50706
rect 59390 50654 59442 50706
rect 59726 50654 59778 50706
rect 60174 50654 60226 50706
rect 64766 50654 64818 50706
rect 65998 50654 66050 50706
rect 69246 50654 69298 50706
rect 73950 50654 74002 50706
rect 80670 50654 80722 50706
rect 97806 50654 97858 50706
rect 51550 50542 51602 50594
rect 53678 50542 53730 50594
rect 55246 50542 55298 50594
rect 56366 50542 56418 50594
rect 56926 50542 56978 50594
rect 57486 50542 57538 50594
rect 58046 50542 58098 50594
rect 61854 50542 61906 50594
rect 71150 50542 71202 50594
rect 74958 50542 75010 50594
rect 75854 50542 75906 50594
rect 79550 50542 79602 50594
rect 83806 50542 83858 50594
rect 91086 50542 91138 50594
rect 92430 50542 92482 50594
rect 93214 50542 93266 50594
rect 93998 50542 94050 50594
rect 95006 50542 95058 50594
rect 50990 50430 51042 50482
rect 52334 50430 52386 50482
rect 52670 50430 52722 50482
rect 54238 50430 54290 50482
rect 62638 50430 62690 50482
rect 65326 50430 65378 50482
rect 70030 50430 70082 50482
rect 71822 50430 71874 50482
rect 77198 50430 77250 50482
rect 85262 50430 85314 50482
rect 85822 50430 85874 50482
rect 87278 50430 87330 50482
rect 88958 50430 89010 50482
rect 89294 50430 89346 50482
rect 89966 50430 90018 50482
rect 90078 50430 90130 50482
rect 91534 50430 91586 50482
rect 91870 50430 91922 50482
rect 94110 50430 94162 50482
rect 95678 50430 95730 50482
rect 51886 50318 51938 50370
rect 52558 50318 52610 50370
rect 53342 50318 53394 50370
rect 53566 50318 53618 50370
rect 54350 50318 54402 50370
rect 54574 50318 54626 50370
rect 57374 50318 57426 50370
rect 65438 50318 65490 50370
rect 65662 50318 65714 50370
rect 66446 50318 66498 50370
rect 69694 50318 69746 50370
rect 69918 50318 69970 50370
rect 70478 50318 70530 50370
rect 75182 50318 75234 50370
rect 76190 50318 76242 50370
rect 89742 50318 89794 50370
rect 90750 50318 90802 50370
rect 90974 50318 91026 50370
rect 91758 50318 91810 50370
rect 93326 50318 93378 50370
rect 94334 50318 94386 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 81278 50150 81330 50202
rect 81382 50150 81434 50202
rect 81486 50150 81538 50202
rect 56702 49982 56754 50034
rect 57598 49982 57650 50034
rect 68350 49982 68402 50034
rect 71934 49982 71986 50034
rect 72158 49982 72210 50034
rect 76414 49982 76466 50034
rect 76862 49982 76914 50034
rect 82350 49982 82402 50034
rect 85038 49982 85090 50034
rect 89406 49982 89458 50034
rect 90190 49982 90242 50034
rect 95566 49982 95618 50034
rect 96126 49982 96178 50034
rect 96350 49982 96402 50034
rect 55582 49870 55634 49922
rect 65550 49870 65602 49922
rect 65662 49870 65714 49922
rect 66334 49870 66386 49922
rect 66894 49870 66946 49922
rect 68910 49870 68962 49922
rect 69358 49870 69410 49922
rect 70590 49870 70642 49922
rect 71486 49870 71538 49922
rect 72270 49870 72322 49922
rect 73390 49870 73442 49922
rect 73726 49870 73778 49922
rect 74286 49870 74338 49922
rect 74622 49870 74674 49922
rect 75182 49870 75234 49922
rect 75518 49870 75570 49922
rect 76078 49870 76130 49922
rect 78318 49870 78370 49922
rect 86494 49870 86546 49922
rect 87614 49870 87666 49922
rect 88398 49870 88450 49922
rect 90302 49870 90354 49922
rect 93326 49870 93378 49922
rect 94782 49870 94834 49922
rect 94894 49870 94946 49922
rect 95454 49870 95506 49922
rect 95790 49870 95842 49922
rect 96462 49870 96514 49922
rect 97358 49870 97410 49922
rect 97470 49870 97522 49922
rect 51886 49758 51938 49810
rect 55358 49758 55410 49810
rect 56478 49758 56530 49810
rect 57486 49758 57538 49810
rect 57822 49758 57874 49810
rect 61854 49758 61906 49810
rect 62526 49758 62578 49810
rect 65326 49758 65378 49810
rect 66446 49758 66498 49810
rect 68014 49758 68066 49810
rect 69694 49758 69746 49810
rect 70366 49758 70418 49810
rect 71262 49758 71314 49810
rect 77534 49758 77586 49810
rect 81790 49758 81842 49810
rect 82238 49758 82290 49810
rect 83022 49758 83074 49810
rect 83582 49758 83634 49810
rect 84366 49758 84418 49810
rect 86382 49758 86434 49810
rect 86718 49758 86770 49810
rect 87502 49758 87554 49810
rect 87838 49758 87890 49810
rect 88286 49758 88338 49810
rect 89294 49758 89346 49810
rect 89630 49758 89682 49810
rect 94110 49758 94162 49810
rect 94558 49758 94610 49810
rect 97134 49758 97186 49810
rect 97918 49758 97970 49810
rect 52558 49646 52610 49698
rect 54686 49646 54738 49698
rect 58158 49646 58210 49698
rect 58606 49646 58658 49698
rect 61294 49646 61346 49698
rect 64654 49646 64706 49698
rect 67454 49646 67506 49698
rect 80446 49646 80498 49698
rect 81342 49646 81394 49698
rect 85486 49646 85538 49698
rect 91198 49646 91250 49698
rect 66334 49534 66386 49586
rect 88398 49534 88450 49586
rect 90190 49534 90242 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 96638 49366 96690 49418
rect 96742 49366 96794 49418
rect 96846 49366 96898 49418
rect 54350 49198 54402 49250
rect 50542 49086 50594 49138
rect 52670 49086 52722 49138
rect 58718 49086 58770 49138
rect 61406 49086 61458 49138
rect 76190 49086 76242 49138
rect 79774 49086 79826 49138
rect 81902 49086 81954 49138
rect 84366 49086 84418 49138
rect 86270 49086 86322 49138
rect 88174 49086 88226 49138
rect 93214 49086 93266 49138
rect 94894 49086 94946 49138
rect 97022 49086 97074 49138
rect 49870 48974 49922 49026
rect 55806 48974 55858 49026
rect 67118 48974 67170 49026
rect 68350 48974 68402 49026
rect 68686 48974 68738 49026
rect 69582 48974 69634 49026
rect 75742 48974 75794 49026
rect 77310 48974 77362 49026
rect 78430 48974 78482 49026
rect 79102 48974 79154 49026
rect 83918 48974 83970 49026
rect 85598 48974 85650 49026
rect 85934 48974 85986 49026
rect 91982 48974 92034 49026
rect 97694 48974 97746 49026
rect 53678 48862 53730 48914
rect 54350 48862 54402 48914
rect 54462 48862 54514 48914
rect 55134 48862 55186 48914
rect 55246 48862 55298 48914
rect 56590 48862 56642 48914
rect 65214 48862 65266 48914
rect 68462 48862 68514 48914
rect 73166 48862 73218 48914
rect 77646 48862 77698 48914
rect 83134 48862 83186 48914
rect 83582 48862 83634 48914
rect 83806 48862 83858 48914
rect 85710 48862 85762 48914
rect 93774 48862 93826 48914
rect 94110 48862 94162 48914
rect 53342 48750 53394 48802
rect 53566 48750 53618 48802
rect 54910 48750 54962 48802
rect 60622 48750 60674 48802
rect 67678 48750 67730 48802
rect 75406 48750 75458 48802
rect 78094 48750 78146 48802
rect 78318 48750 78370 48802
rect 82350 48750 82402 48802
rect 82798 48750 82850 48802
rect 83022 48750 83074 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 81278 48582 81330 48634
rect 81382 48582 81434 48634
rect 81486 48582 81538 48634
rect 53342 48414 53394 48466
rect 53902 48414 53954 48466
rect 57598 48414 57650 48466
rect 58606 48414 58658 48466
rect 61854 48414 61906 48466
rect 62638 48414 62690 48466
rect 63198 48414 63250 48466
rect 64206 48414 64258 48466
rect 67342 48414 67394 48466
rect 68014 48414 68066 48466
rect 72046 48414 72098 48466
rect 78318 48414 78370 48466
rect 92654 48414 92706 48466
rect 97918 48414 97970 48466
rect 50542 48302 50594 48354
rect 53454 48302 53506 48354
rect 54126 48302 54178 48354
rect 54910 48302 54962 48354
rect 55022 48302 55074 48354
rect 56478 48302 56530 48354
rect 57374 48302 57426 48354
rect 58270 48302 58322 48354
rect 58382 48302 58434 48354
rect 59166 48302 59218 48354
rect 60734 48302 60786 48354
rect 62526 48302 62578 48354
rect 62862 48302 62914 48354
rect 63422 48302 63474 48354
rect 63534 48302 63586 48354
rect 65550 48302 65602 48354
rect 66334 48302 66386 48354
rect 69470 48302 69522 48354
rect 72270 48302 72322 48354
rect 72382 48302 72434 48354
rect 78766 48302 78818 48354
rect 82350 48302 82402 48354
rect 87166 48302 87218 48354
rect 90078 48302 90130 48354
rect 92878 48302 92930 48354
rect 92990 48302 93042 48354
rect 97358 48302 97410 48354
rect 97470 48302 97522 48354
rect 49870 48190 49922 48242
rect 53118 48190 53170 48242
rect 54238 48190 54290 48242
rect 56254 48190 56306 48242
rect 56590 48190 56642 48242
rect 57710 48190 57762 48242
rect 58942 48190 58994 48242
rect 59278 48190 59330 48242
rect 60622 48190 60674 48242
rect 60958 48190 61010 48242
rect 61966 48190 62018 48242
rect 64318 48190 64370 48242
rect 65326 48190 65378 48242
rect 65662 48190 65714 48242
rect 66110 48190 66162 48242
rect 66446 48190 66498 48242
rect 67902 48190 67954 48242
rect 68238 48190 68290 48242
rect 68686 48190 68738 48242
rect 76750 48190 76802 48242
rect 77646 48190 77698 48242
rect 78094 48190 78146 48242
rect 79550 48190 79602 48242
rect 80446 48190 80498 48242
rect 81678 48190 81730 48242
rect 87950 48190 88002 48242
rect 89294 48190 89346 48242
rect 93662 48190 93714 48242
rect 52670 48078 52722 48130
rect 55470 48078 55522 48130
rect 59726 48078 59778 48130
rect 66894 48078 66946 48130
rect 71598 48078 71650 48130
rect 73278 48078 73330 48130
rect 73838 48078 73890 48130
rect 75966 48078 76018 48130
rect 77310 48078 77362 48130
rect 84478 48078 84530 48130
rect 85038 48078 85090 48130
rect 88622 48078 88674 48130
rect 92206 48078 92258 48130
rect 94334 48078 94386 48130
rect 96462 48078 96514 48130
rect 54910 47966 54962 48018
rect 61854 47966 61906 48018
rect 64206 47966 64258 48018
rect 97358 47966 97410 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 96638 47798 96690 47850
rect 96742 47798 96794 47850
rect 96846 47798 96898 47850
rect 50094 47518 50146 47570
rect 52222 47518 52274 47570
rect 55806 47518 55858 47570
rect 59950 47518 60002 47570
rect 60622 47518 60674 47570
rect 62078 47518 62130 47570
rect 62862 47518 62914 47570
rect 67006 47518 67058 47570
rect 67790 47518 67842 47570
rect 70814 47518 70866 47570
rect 75854 47518 75906 47570
rect 76414 47518 76466 47570
rect 78654 47518 78706 47570
rect 81006 47518 81058 47570
rect 82238 47518 82290 47570
rect 83470 47518 83522 47570
rect 84142 47518 84194 47570
rect 84478 47518 84530 47570
rect 89966 47518 90018 47570
rect 92094 47518 92146 47570
rect 94782 47518 94834 47570
rect 97246 47518 97298 47570
rect 49422 47406 49474 47458
rect 54910 47406 54962 47458
rect 61742 47406 61794 47458
rect 65774 47406 65826 47458
rect 66558 47406 66610 47458
rect 69582 47406 69634 47458
rect 72158 47406 72210 47458
rect 73054 47418 73106 47470
rect 77198 47406 77250 47458
rect 85598 47406 85650 47458
rect 86494 47406 86546 47458
rect 86942 47406 86994 47458
rect 87726 47406 87778 47458
rect 88174 47406 88226 47458
rect 89294 47406 89346 47458
rect 96126 47406 96178 47458
rect 96462 47406 96514 47458
rect 61406 47294 61458 47346
rect 61518 47294 61570 47346
rect 64990 47294 65042 47346
rect 68462 47294 68514 47346
rect 68574 47294 68626 47346
rect 69470 47294 69522 47346
rect 70030 47294 70082 47346
rect 70366 47294 70418 47346
rect 72270 47294 72322 47346
rect 73726 47294 73778 47346
rect 78206 47294 78258 47346
rect 88622 47294 88674 47346
rect 93214 47294 93266 47346
rect 93550 47294 93602 47346
rect 94334 47294 94386 47346
rect 95230 47294 95282 47346
rect 96238 47294 96290 47346
rect 52670 47182 52722 47234
rect 59502 47182 59554 47234
rect 66222 47182 66274 47234
rect 66446 47182 66498 47234
rect 68238 47182 68290 47234
rect 69246 47182 69298 47234
rect 70254 47182 70306 47234
rect 71262 47182 71314 47234
rect 72494 47182 72546 47234
rect 77646 47182 77698 47234
rect 87614 47182 87666 47234
rect 93998 47182 94050 47234
rect 94222 47182 94274 47234
rect 96798 47182 96850 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 81278 47014 81330 47066
rect 81382 47014 81434 47066
rect 81486 47014 81538 47066
rect 53342 46846 53394 46898
rect 53566 46846 53618 46898
rect 54238 46846 54290 46898
rect 55246 46846 55298 46898
rect 55694 46846 55746 46898
rect 56030 46846 56082 46898
rect 57486 46846 57538 46898
rect 66222 46846 66274 46898
rect 70590 46846 70642 46898
rect 71934 46846 71986 46898
rect 72718 46846 72770 46898
rect 73278 46846 73330 46898
rect 73950 46846 74002 46898
rect 75630 46846 75682 46898
rect 75854 46846 75906 46898
rect 76414 46846 76466 46898
rect 77534 46846 77586 46898
rect 77982 46846 78034 46898
rect 82462 46846 82514 46898
rect 85150 46846 85202 46898
rect 93214 46846 93266 46898
rect 93438 46846 93490 46898
rect 93774 46846 93826 46898
rect 95118 46846 95170 46898
rect 95678 46846 95730 46898
rect 96014 46846 96066 46898
rect 96574 46846 96626 46898
rect 53678 46734 53730 46786
rect 62190 46734 62242 46786
rect 65550 46734 65602 46786
rect 65662 46734 65714 46786
rect 73838 46734 73890 46786
rect 75070 46734 75122 46786
rect 75518 46734 75570 46786
rect 76302 46734 76354 46786
rect 87726 46734 87778 46786
rect 93102 46734 93154 46786
rect 61518 46622 61570 46674
rect 66894 46622 66946 46674
rect 82238 46622 82290 46674
rect 88398 46622 88450 46674
rect 89630 46622 89682 46674
rect 52446 46510 52498 46562
rect 52894 46510 52946 46562
rect 54798 46510 54850 46562
rect 60958 46510 61010 46562
rect 64318 46510 64370 46562
rect 67566 46510 67618 46562
rect 69694 46510 69746 46562
rect 70142 46510 70194 46562
rect 76974 46510 77026 46562
rect 81678 46510 81730 46562
rect 85598 46510 85650 46562
rect 90414 46510 90466 46562
rect 92542 46510 92594 46562
rect 94334 46510 94386 46562
rect 94782 46510 94834 46562
rect 54462 46398 54514 46450
rect 54798 46398 54850 46450
rect 55470 46398 55522 46450
rect 56030 46398 56082 46450
rect 65550 46398 65602 46450
rect 73950 46398 74002 46450
rect 76414 46398 76466 46450
rect 94782 46398 94834 46450
rect 95678 46398 95730 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 64990 46062 65042 46114
rect 94334 46062 94386 46114
rect 95342 46062 95394 46114
rect 56142 45950 56194 46002
rect 58270 45950 58322 46002
rect 62190 45950 62242 46002
rect 64318 45950 64370 46002
rect 75294 45950 75346 46002
rect 76078 45950 76130 46002
rect 83918 45950 83970 46002
rect 89070 45950 89122 46002
rect 91310 45950 91362 46002
rect 92430 45950 92482 46002
rect 94110 45950 94162 46002
rect 94670 45950 94722 46002
rect 95118 45950 95170 46002
rect 55470 45838 55522 45890
rect 61518 45838 61570 45890
rect 65102 45838 65154 45890
rect 68126 45838 68178 45890
rect 68462 45838 68514 45890
rect 81342 45838 81394 45890
rect 82238 45838 82290 45890
rect 82574 45838 82626 45890
rect 85710 45838 85762 45890
rect 89742 45838 89794 45890
rect 90078 45838 90130 45890
rect 90526 45838 90578 45890
rect 90862 45838 90914 45890
rect 51214 45726 51266 45778
rect 64990 45726 65042 45778
rect 68350 45726 68402 45778
rect 79102 45726 79154 45778
rect 80670 45726 80722 45778
rect 82798 45726 82850 45778
rect 83134 45726 83186 45778
rect 84478 45726 84530 45778
rect 85934 45726 85986 45778
rect 86270 45726 86322 45778
rect 89854 45726 89906 45778
rect 90750 45726 90802 45778
rect 50878 45614 50930 45666
rect 58718 45614 58770 45666
rect 70142 45614 70194 45666
rect 77310 45614 77362 45666
rect 78766 45614 78818 45666
rect 81566 45614 81618 45666
rect 85374 45614 85426 45666
rect 91982 45614 92034 45666
rect 93102 45614 93154 45666
rect 93550 45614 93602 45666
rect 95566 45614 95618 45666
rect 95902 45614 95954 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 70926 45278 70978 45330
rect 71374 45278 71426 45330
rect 74734 45278 74786 45330
rect 75070 45278 75122 45330
rect 50766 45166 50818 45218
rect 56254 45166 56306 45218
rect 63534 45166 63586 45218
rect 67678 45166 67730 45218
rect 75630 45166 75682 45218
rect 77086 45166 77138 45218
rect 78430 45166 78482 45218
rect 82126 45166 82178 45218
rect 91982 45166 92034 45218
rect 96126 45166 96178 45218
rect 50094 45054 50146 45106
rect 56590 45054 56642 45106
rect 64206 45054 64258 45106
rect 67006 45054 67058 45106
rect 75966 45054 76018 45106
rect 76750 45054 76802 45106
rect 77758 45054 77810 45106
rect 81342 45054 81394 45106
rect 84926 45054 84978 45106
rect 91422 45054 91474 45106
rect 95790 45054 95842 45106
rect 52894 44942 52946 44994
rect 53454 44942 53506 44994
rect 61406 44942 61458 44994
rect 69806 44942 69858 44994
rect 70366 44942 70418 44994
rect 80558 44942 80610 44994
rect 84254 44942 84306 44994
rect 85598 44942 85650 44994
rect 87726 44942 87778 44994
rect 88174 44942 88226 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 77422 44494 77474 44546
rect 93326 44494 93378 44546
rect 93998 44494 94050 44546
rect 51886 44382 51938 44434
rect 56030 44382 56082 44434
rect 58158 44382 58210 44434
rect 58606 44382 58658 44434
rect 59278 44382 59330 44434
rect 61854 44382 61906 44434
rect 72382 44382 72434 44434
rect 74398 44382 74450 44434
rect 76526 44382 76578 44434
rect 77758 44382 77810 44434
rect 80670 44382 80722 44434
rect 93102 44382 93154 44434
rect 93998 44382 94050 44434
rect 94894 44382 94946 44434
rect 97022 44382 97074 44434
rect 49086 44270 49138 44322
rect 55358 44270 55410 44322
rect 62526 44270 62578 44322
rect 67230 44270 67282 44322
rect 69470 44270 69522 44322
rect 73726 44270 73778 44322
rect 83918 44270 83970 44322
rect 85374 44270 85426 44322
rect 91310 44270 91362 44322
rect 91982 44270 92034 44322
rect 93550 44270 93602 44322
rect 97694 44270 97746 44322
rect 49758 44158 49810 44210
rect 66334 44158 66386 44210
rect 70254 44158 70306 44210
rect 77982 44158 78034 44210
rect 78542 44158 78594 44210
rect 85598 44158 85650 44210
rect 91198 44158 91250 44210
rect 52334 44046 52386 44098
rect 62750 44046 62802 44098
rect 72830 44046 72882 44098
rect 90638 44046 90690 44098
rect 92318 44046 92370 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 48750 43710 48802 43762
rect 63422 43710 63474 43762
rect 70254 43710 70306 43762
rect 76302 43710 76354 43762
rect 50766 43598 50818 43650
rect 51662 43598 51714 43650
rect 52222 43598 52274 43650
rect 52782 43598 52834 43650
rect 54350 43598 54402 43650
rect 55022 43598 55074 43650
rect 56702 43598 56754 43650
rect 57598 43598 57650 43650
rect 58494 43598 58546 43650
rect 59838 43598 59890 43650
rect 64430 43598 64482 43650
rect 71486 43598 71538 43650
rect 72046 43598 72098 43650
rect 72718 43598 72770 43650
rect 75294 43598 75346 43650
rect 77870 43598 77922 43650
rect 95566 43598 95618 43650
rect 97134 43598 97186 43650
rect 48526 43486 48578 43538
rect 49758 43486 49810 43538
rect 50878 43486 50930 43538
rect 53790 43486 53842 43538
rect 55358 43486 55410 43538
rect 58718 43486 58770 43538
rect 60174 43486 60226 43538
rect 64542 43486 64594 43538
rect 65774 43486 65826 43538
rect 70030 43486 70082 43538
rect 70926 43486 70978 43538
rect 71262 43486 71314 43538
rect 74622 43486 74674 43538
rect 75182 43486 75234 43538
rect 75966 43486 76018 43538
rect 77198 43486 77250 43538
rect 92654 43486 92706 43538
rect 50094 43374 50146 43426
rect 51998 43374 52050 43426
rect 53342 43374 53394 43426
rect 59278 43374 59330 43426
rect 65326 43374 65378 43426
rect 69358 43374 69410 43426
rect 79998 43374 80050 43426
rect 84702 43374 84754 43426
rect 89742 43374 89794 43426
rect 90078 43374 90130 43426
rect 57934 43262 57986 43314
rect 63758 43262 63810 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 77422 42926 77474 42978
rect 77758 42926 77810 42978
rect 52670 42814 52722 42866
rect 53454 42814 53506 42866
rect 54798 42814 54850 42866
rect 56926 42814 56978 42866
rect 60398 42814 60450 42866
rect 62526 42814 62578 42866
rect 63870 42814 63922 42866
rect 65998 42814 66050 42866
rect 68574 42814 68626 42866
rect 72270 42814 72322 42866
rect 79214 42814 79266 42866
rect 87502 42814 87554 42866
rect 94334 42814 94386 42866
rect 94894 42814 94946 42866
rect 49758 42702 49810 42754
rect 54126 42702 54178 42754
rect 57598 42702 57650 42754
rect 63086 42702 63138 42754
rect 69358 42702 69410 42754
rect 75742 42702 75794 42754
rect 81790 42702 81842 42754
rect 86158 42702 86210 42754
rect 89742 42702 89794 42754
rect 93214 42702 93266 42754
rect 97694 42702 97746 42754
rect 50542 42590 50594 42642
rect 58270 42590 58322 42642
rect 77982 42590 78034 42642
rect 78542 42590 78594 42642
rect 85262 42590 85314 42642
rect 86382 42590 86434 42642
rect 86942 42590 86994 42642
rect 89966 42590 90018 42642
rect 90526 42590 90578 42642
rect 97022 42590 97074 42642
rect 61294 42478 61346 42530
rect 62078 42478 62130 42530
rect 66446 42478 66498 42530
rect 75182 42478 75234 42530
rect 76190 42478 76242 42530
rect 82014 42478 82066 42530
rect 85822 42478 85874 42530
rect 88286 42478 88338 42530
rect 88734 42478 88786 42530
rect 89406 42478 89458 42530
rect 92430 42478 92482 42530
rect 93550 42478 93602 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 54798 42142 54850 42194
rect 71710 42142 71762 42194
rect 77758 42142 77810 42194
rect 97246 42142 97298 42194
rect 54126 42030 54178 42082
rect 56590 42030 56642 42082
rect 60734 42030 60786 42082
rect 64318 42030 64370 42082
rect 65438 42030 65490 42082
rect 65774 42030 65826 42082
rect 70814 42030 70866 42082
rect 82126 42030 82178 42082
rect 95342 42030 95394 42082
rect 49646 41918 49698 41970
rect 54238 41918 54290 41970
rect 55470 41918 55522 41970
rect 56478 41918 56530 41970
rect 62078 41918 62130 41970
rect 64430 41918 64482 41970
rect 66334 41918 66386 41970
rect 70926 41918 70978 41970
rect 73278 41918 73330 41970
rect 73950 41918 74002 41970
rect 81342 41918 81394 41970
rect 84926 41918 84978 41970
rect 88174 41918 88226 41970
rect 89294 41918 89346 41970
rect 95230 41918 95282 41970
rect 96350 41918 96402 41970
rect 97470 41918 97522 41970
rect 98030 41918 98082 41970
rect 50318 41806 50370 41858
rect 52446 41806 52498 41858
rect 53454 41806 53506 41858
rect 63422 41806 63474 41858
rect 67118 41806 67170 41858
rect 69246 41806 69298 41858
rect 72158 41806 72210 41858
rect 74734 41806 74786 41858
rect 76862 41806 76914 41858
rect 77310 41806 77362 41858
rect 78206 41806 78258 41858
rect 84254 41806 84306 41858
rect 85598 41806 85650 41858
rect 87726 41806 87778 41858
rect 94334 41806 94386 41858
rect 53118 41694 53170 41746
rect 55806 41694 55858 41746
rect 63758 41694 63810 41746
rect 69918 41694 69970 41746
rect 70254 41694 70306 41746
rect 96014 41694 96066 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 51774 41358 51826 41410
rect 53230 41358 53282 41410
rect 53790 41358 53842 41410
rect 58942 41358 58994 41410
rect 82126 41358 82178 41410
rect 90302 41358 90354 41410
rect 53342 41246 53394 41298
rect 53790 41246 53842 41298
rect 54238 41246 54290 41298
rect 55134 41246 55186 41298
rect 56590 41246 56642 41298
rect 56926 41246 56978 41298
rect 62190 41246 62242 41298
rect 64318 41246 64370 41298
rect 65550 41246 65602 41298
rect 68686 41246 68738 41298
rect 69470 41246 69522 41298
rect 70366 41246 70418 41298
rect 70814 41246 70866 41298
rect 72270 41246 72322 41298
rect 72718 41246 72770 41298
rect 75854 41246 75906 41298
rect 84254 41246 84306 41298
rect 86718 41246 86770 41298
rect 93214 41246 93266 41298
rect 95342 41246 95394 41298
rect 50766 41134 50818 41186
rect 52558 41134 52610 41186
rect 57710 41134 57762 41186
rect 58606 41134 58658 41186
rect 59726 41134 59778 41186
rect 60286 41134 60338 41186
rect 64990 41134 65042 41186
rect 65998 41134 66050 41186
rect 67678 41134 67730 41186
rect 71822 41134 71874 41186
rect 73838 41134 73890 41186
rect 77534 41134 77586 41186
rect 82462 41134 82514 41186
rect 85822 41134 85874 41186
rect 89630 41134 89682 41186
rect 90638 41134 90690 41186
rect 91310 41134 91362 41186
rect 96126 41134 96178 41186
rect 97134 41134 97186 41186
rect 97582 41134 97634 41186
rect 49534 41022 49586 41074
rect 49870 41022 49922 41074
rect 50430 41022 50482 41074
rect 51438 41022 51490 41074
rect 52334 41022 52386 41074
rect 54686 41022 54738 41074
rect 57934 41022 57986 41074
rect 59502 41022 59554 41074
rect 67342 41022 67394 41074
rect 74062 41022 74114 41074
rect 74622 41022 74674 41074
rect 77310 41022 77362 41074
rect 78990 41022 79042 41074
rect 81566 41022 81618 41074
rect 82686 41022 82738 41074
rect 83246 41022 83298 41074
rect 85598 41022 85650 41074
rect 88846 41022 88898 41074
rect 91198 41022 91250 41074
rect 92430 41022 92482 41074
rect 96798 41022 96850 41074
rect 97918 41022 97970 41074
rect 69918 40910 69970 40962
rect 73502 40910 73554 40962
rect 75294 40910 75346 40962
rect 76302 40910 76354 40962
rect 79326 40910 79378 40962
rect 83806 40910 83858 40962
rect 92094 40910 92146 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 62190 40574 62242 40626
rect 62750 40574 62802 40626
rect 64542 40574 64594 40626
rect 70702 40574 70754 40626
rect 71262 40574 71314 40626
rect 72270 40574 72322 40626
rect 74174 40574 74226 40626
rect 74622 40574 74674 40626
rect 89294 40574 89346 40626
rect 98030 40574 98082 40626
rect 53342 40462 53394 40514
rect 59614 40462 59666 40514
rect 63534 40462 63586 40514
rect 63982 40462 64034 40514
rect 73390 40462 73442 40514
rect 88174 40462 88226 40514
rect 96126 40462 96178 40514
rect 97246 40462 97298 40514
rect 55582 40350 55634 40402
rect 56030 40350 56082 40402
rect 58158 40350 58210 40402
rect 58942 40350 58994 40402
rect 65326 40350 65378 40402
rect 67454 40350 67506 40402
rect 73614 40350 73666 40402
rect 80446 40350 80498 40402
rect 81230 40350 81282 40402
rect 82686 40350 82738 40402
rect 83918 40350 83970 40402
rect 89518 40350 89570 40402
rect 95678 40350 95730 40402
rect 97470 40350 97522 40402
rect 61742 40238 61794 40290
rect 64206 40238 64258 40290
rect 68126 40238 68178 40290
rect 70254 40238 70306 40290
rect 71710 40238 71762 40290
rect 77758 40238 77810 40290
rect 90862 40238 90914 40290
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 64990 39678 65042 39730
rect 70702 39678 70754 39730
rect 72718 39678 72770 39730
rect 74846 39678 74898 39730
rect 75854 39678 75906 39730
rect 77198 39678 77250 39730
rect 79214 39678 79266 39730
rect 81342 39678 81394 39730
rect 85150 39678 85202 39730
rect 87950 39678 88002 39730
rect 93326 39678 93378 39730
rect 94894 39678 94946 39730
rect 97022 39678 97074 39730
rect 53454 39566 53506 39618
rect 61742 39566 61794 39618
rect 62302 39566 62354 39618
rect 69694 39566 69746 39618
rect 70254 39566 70306 39618
rect 72046 39566 72098 39618
rect 75406 39566 75458 39618
rect 76414 39566 76466 39618
rect 78430 39566 78482 39618
rect 82350 39566 82402 39618
rect 83246 39566 83298 39618
rect 83582 39566 83634 39618
rect 84142 39566 84194 39618
rect 90862 39566 90914 39618
rect 93886 39566 93938 39618
rect 97806 39566 97858 39618
rect 51102 39454 51154 39506
rect 51438 39454 51490 39506
rect 55806 39454 55858 39506
rect 59950 39454 60002 39506
rect 68238 39454 68290 39506
rect 68574 39454 68626 39506
rect 84366 39454 84418 39506
rect 90078 39454 90130 39506
rect 50542 39342 50594 39394
rect 55470 39342 55522 39394
rect 59614 39342 59666 39394
rect 61294 39342 61346 39394
rect 77870 39342 77922 39394
rect 82574 39342 82626 39394
rect 94222 39342 94274 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 62190 39006 62242 39058
rect 69694 39006 69746 39058
rect 71374 39006 71426 39058
rect 78990 39006 79042 39058
rect 81342 39006 81394 39058
rect 85822 39006 85874 39058
rect 88510 39006 88562 39058
rect 89630 39006 89682 39058
rect 94558 39006 94610 39058
rect 96350 39006 96402 39058
rect 97134 39006 97186 39058
rect 97582 39006 97634 39058
rect 50318 38894 50370 38946
rect 52222 38894 52274 38946
rect 53006 38894 53058 38946
rect 54574 38894 54626 38946
rect 59390 38894 59442 38946
rect 63086 38894 63138 38946
rect 63982 38894 64034 38946
rect 70814 38894 70866 38946
rect 74846 38894 74898 38946
rect 76190 38894 76242 38946
rect 80110 38894 80162 38946
rect 83246 38894 83298 38946
rect 90526 38894 90578 38946
rect 91870 38894 91922 38946
rect 95454 38894 95506 38946
rect 50654 38782 50706 38834
rect 51326 38782 51378 38834
rect 52446 38782 52498 38834
rect 53790 38782 53842 38834
rect 58718 38782 58770 38834
rect 62526 38782 62578 38834
rect 63198 38782 63250 38834
rect 64206 38782 64258 38834
rect 65550 38782 65602 38834
rect 70030 38782 70082 38834
rect 70702 38782 70754 38834
rect 74622 38782 74674 38834
rect 75518 38782 75570 38834
rect 79998 38782 80050 38834
rect 82574 38782 82626 38834
rect 89406 38782 89458 38834
rect 90190 38782 90242 38834
rect 91198 38782 91250 38834
rect 95230 38782 95282 38834
rect 96014 38782 96066 38834
rect 56702 38670 56754 38722
rect 61518 38670 61570 38722
rect 66222 38670 66274 38722
rect 68350 38670 68402 38722
rect 71822 38670 71874 38722
rect 78318 38670 78370 38722
rect 79326 38670 79378 38722
rect 85374 38670 85426 38722
rect 93998 38670 94050 38722
rect 98030 38670 98082 38722
rect 51662 38558 51714 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 56366 38222 56418 38274
rect 56702 38222 56754 38274
rect 74846 38222 74898 38274
rect 75182 38222 75234 38274
rect 50542 38110 50594 38162
rect 52670 38110 52722 38162
rect 53454 38110 53506 38162
rect 53790 38110 53842 38162
rect 61518 38110 61570 38162
rect 62862 38110 62914 38162
rect 64990 38110 65042 38162
rect 65550 38110 65602 38162
rect 69246 38110 69298 38162
rect 69694 38110 69746 38162
rect 76526 38110 76578 38162
rect 78990 38110 79042 38162
rect 84254 38110 84306 38162
rect 85150 38110 85202 38162
rect 93326 38110 93378 38162
rect 97582 38110 97634 38162
rect 98030 38110 98082 38162
rect 48974 37998 49026 38050
rect 49758 37998 49810 38050
rect 57374 37998 57426 38050
rect 62190 37998 62242 38050
rect 67566 37998 67618 38050
rect 68350 37998 68402 38050
rect 75854 37998 75906 38050
rect 77310 37998 77362 38050
rect 77870 37998 77922 38050
rect 78542 37998 78594 38050
rect 81454 37998 81506 38050
rect 89182 37998 89234 38050
rect 90974 37998 91026 38050
rect 91646 37998 91698 38050
rect 94670 37998 94722 38050
rect 1822 37886 1874 37938
rect 2158 37886 2210 37938
rect 57262 37886 57314 37938
rect 66222 37886 66274 37938
rect 66558 37886 66610 37938
rect 67230 37886 67282 37938
rect 68238 37886 68290 37938
rect 75966 37886 76018 37938
rect 82126 37886 82178 37938
rect 90862 37886 90914 37938
rect 93774 37886 93826 37938
rect 94110 37886 94162 37938
rect 95454 37886 95506 37938
rect 49198 37774 49250 37826
rect 55694 37774 55746 37826
rect 58046 37774 58098 37826
rect 88510 37774 88562 37826
rect 89406 37774 89458 37826
rect 89854 37774 89906 37826
rect 91982 37774 92034 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 1822 37438 1874 37490
rect 52894 37438 52946 37490
rect 59390 37438 59442 37490
rect 59838 37438 59890 37490
rect 63422 37438 63474 37490
rect 65326 37438 65378 37490
rect 65774 37438 65826 37490
rect 74174 37438 74226 37490
rect 75294 37438 75346 37490
rect 77086 37438 77138 37490
rect 81902 37438 81954 37490
rect 93886 37438 93938 37490
rect 94222 37438 94274 37490
rect 96350 37438 96402 37490
rect 50318 37326 50370 37378
rect 56702 37326 56754 37378
rect 58830 37326 58882 37378
rect 64318 37326 64370 37378
rect 75854 37326 75906 37378
rect 76414 37326 76466 37378
rect 77870 37326 77922 37378
rect 83806 37326 83858 37378
rect 91422 37326 91474 37378
rect 92766 37326 92818 37378
rect 93102 37326 93154 37378
rect 95342 37326 95394 37378
rect 49646 37214 49698 37266
rect 56478 37214 56530 37266
rect 57710 37214 57762 37266
rect 58718 37214 58770 37266
rect 64430 37214 64482 37266
rect 66782 37214 66834 37266
rect 75630 37214 75682 37266
rect 82238 37214 82290 37266
rect 82910 37214 82962 37266
rect 83246 37214 83298 37266
rect 83918 37214 83970 37266
rect 92206 37214 92258 37266
rect 95454 37214 95506 37266
rect 96014 37214 96066 37266
rect 52446 37102 52498 37154
rect 67454 37102 67506 37154
rect 69582 37102 69634 37154
rect 70142 37102 70194 37154
rect 74622 37102 74674 37154
rect 77422 37102 77474 37154
rect 84590 37102 84642 37154
rect 89294 37102 89346 37154
rect 97134 37102 97186 37154
rect 58046 36990 58098 37042
rect 63758 36990 63810 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 51102 36654 51154 36706
rect 51438 36654 51490 36706
rect 64878 36654 64930 36706
rect 65438 36654 65490 36706
rect 69806 36654 69858 36706
rect 95230 36654 95282 36706
rect 95566 36654 95618 36706
rect 53790 36542 53842 36594
rect 56814 36542 56866 36594
rect 58942 36542 58994 36594
rect 61518 36542 61570 36594
rect 64990 36542 65042 36594
rect 65438 36542 65490 36594
rect 71150 36542 71202 36594
rect 73390 36542 73442 36594
rect 74286 36542 74338 36594
rect 77198 36542 77250 36594
rect 77646 36542 77698 36594
rect 82574 36542 82626 36594
rect 87054 36542 87106 36594
rect 89518 36542 89570 36594
rect 91646 36542 91698 36594
rect 93214 36542 93266 36594
rect 96910 36542 96962 36594
rect 52222 36430 52274 36482
rect 53342 36430 53394 36482
rect 56142 36430 56194 36482
rect 70590 36430 70642 36482
rect 73838 36430 73890 36482
rect 74958 36430 75010 36482
rect 75406 36430 75458 36482
rect 76078 36430 76130 36482
rect 92430 36430 92482 36482
rect 93774 36430 93826 36482
rect 94334 36430 94386 36482
rect 52110 36318 52162 36370
rect 59502 36318 59554 36370
rect 68014 36318 68066 36370
rect 68350 36318 68402 36370
rect 69470 36318 69522 36370
rect 70366 36318 70418 36370
rect 71598 36318 71650 36370
rect 76414 36318 76466 36370
rect 95790 36318 95842 36370
rect 96238 36318 96290 36370
rect 54238 36206 54290 36258
rect 59838 36206 59890 36258
rect 60286 36206 60338 36258
rect 94558 36206 94610 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 55246 35870 55298 35922
rect 56702 35870 56754 35922
rect 59054 35870 59106 35922
rect 59726 35870 59778 35922
rect 61070 35870 61122 35922
rect 64542 35870 64594 35922
rect 74062 35870 74114 35922
rect 77310 35870 77362 35922
rect 81230 35870 81282 35922
rect 81678 35870 81730 35922
rect 82462 35870 82514 35922
rect 84478 35870 84530 35922
rect 84926 35870 84978 35922
rect 89406 35870 89458 35922
rect 54126 35758 54178 35810
rect 54462 35758 54514 35810
rect 58046 35758 58098 35810
rect 58494 35758 58546 35810
rect 60622 35758 60674 35810
rect 61966 35758 62018 35810
rect 62526 35758 62578 35810
rect 71710 35758 71762 35810
rect 74958 35758 75010 35810
rect 76526 35758 76578 35810
rect 83358 35758 83410 35810
rect 86158 35758 86210 35810
rect 86718 35758 86770 35810
rect 87614 35758 87666 35810
rect 88510 35758 88562 35810
rect 89966 35758 90018 35810
rect 90302 35758 90354 35810
rect 97134 35758 97186 35810
rect 49982 35646 50034 35698
rect 60286 35646 60338 35698
rect 62750 35646 62802 35698
rect 63086 35646 63138 35698
rect 71934 35646 71986 35698
rect 74734 35646 74786 35698
rect 76750 35646 76802 35698
rect 83134 35646 83186 35698
rect 87838 35646 87890 35698
rect 89742 35646 89794 35698
rect 96462 35646 96514 35698
rect 50766 35534 50818 35586
rect 52894 35534 52946 35586
rect 63646 35534 63698 35586
rect 66670 35534 66722 35586
rect 72606 35534 72658 35586
rect 73502 35534 73554 35586
rect 75854 35534 75906 35586
rect 94446 35534 94498 35586
rect 53566 35422 53618 35474
rect 53902 35422 53954 35474
rect 58718 35422 58770 35474
rect 75518 35422 75570 35474
rect 84478 35422 84530 35474
rect 85262 35422 85314 35474
rect 85598 35422 85650 35474
rect 85934 35422 85986 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 71822 35086 71874 35138
rect 52670 34974 52722 35026
rect 53454 34974 53506 35026
rect 57374 34974 57426 35026
rect 62190 34974 62242 35026
rect 64318 34974 64370 35026
rect 66670 34974 66722 35026
rect 74398 34974 74450 35026
rect 76526 34974 76578 35026
rect 81678 34974 81730 35026
rect 88174 34974 88226 35026
rect 88622 34974 88674 35026
rect 90302 34974 90354 35026
rect 97246 34974 97298 35026
rect 49870 34862 49922 34914
rect 56814 34862 56866 34914
rect 61406 34862 61458 34914
rect 65326 34862 65378 34914
rect 66110 34862 66162 34914
rect 67678 34862 67730 34914
rect 68462 34862 68514 34914
rect 69694 34862 69746 34914
rect 72158 34862 72210 34914
rect 73726 34862 73778 34914
rect 77310 34862 77362 34914
rect 78766 34862 78818 34914
rect 82686 34862 82738 34914
rect 84254 34862 84306 34914
rect 85262 34862 85314 34914
rect 90974 34862 91026 34914
rect 91646 34862 91698 34914
rect 94446 34862 94498 34914
rect 50542 34750 50594 34802
rect 54350 34750 54402 34802
rect 54686 34750 54738 34802
rect 65886 34750 65938 34802
rect 68238 34750 68290 34802
rect 71150 34750 71202 34802
rect 72382 34750 72434 34802
rect 72718 34750 72770 34802
rect 79550 34750 79602 34802
rect 82910 34750 82962 34802
rect 83246 34750 83298 34802
rect 84478 34750 84530 34802
rect 86046 34750 86098 34802
rect 90862 34750 90914 34802
rect 95118 34750 95170 34802
rect 53790 34638 53842 34690
rect 64990 34638 65042 34690
rect 67342 34638 67394 34690
rect 69358 34638 69410 34690
rect 70814 34638 70866 34690
rect 82350 34638 82402 34690
rect 89854 34638 89906 34690
rect 91982 34638 92034 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 50990 34302 51042 34354
rect 64542 34302 64594 34354
rect 66222 34302 66274 34354
rect 73502 34302 73554 34354
rect 75294 34302 75346 34354
rect 79550 34302 79602 34354
rect 93662 34302 93714 34354
rect 94558 34302 94610 34354
rect 95230 34302 95282 34354
rect 97134 34302 97186 34354
rect 51326 34190 51378 34242
rect 53006 34190 53058 34242
rect 59614 34190 59666 34242
rect 65438 34190 65490 34242
rect 65774 34190 65826 34242
rect 70142 34190 70194 34242
rect 74398 34190 74450 34242
rect 79886 34190 79938 34242
rect 87950 34190 88002 34242
rect 88174 34190 88226 34242
rect 92766 34190 92818 34242
rect 93102 34190 93154 34242
rect 95790 34190 95842 34242
rect 96126 34190 96178 34242
rect 52334 34078 52386 34130
rect 53118 34078 53170 34130
rect 53902 34078 53954 34130
rect 60286 34078 60338 34130
rect 60958 34078 61010 34130
rect 67230 34078 67282 34130
rect 73838 34078 73890 34130
rect 74622 34078 74674 34130
rect 78766 34078 78818 34130
rect 86606 34078 86658 34130
rect 89406 34078 89458 34130
rect 94334 34078 94386 34130
rect 95566 34078 95618 34130
rect 54574 33966 54626 34018
rect 56702 33966 56754 34018
rect 57486 33966 57538 34018
rect 61742 33966 61794 34018
rect 63870 33966 63922 34018
rect 75966 33966 76018 34018
rect 78094 33966 78146 34018
rect 82462 33966 82514 34018
rect 87614 33966 87666 34018
rect 90078 33966 90130 34018
rect 92206 33966 92258 34018
rect 51998 33854 52050 33906
rect 87278 33854 87330 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 72830 33518 72882 33570
rect 73502 33518 73554 33570
rect 82126 33518 82178 33570
rect 53454 33406 53506 33458
rect 53790 33406 53842 33458
rect 57374 33406 57426 33458
rect 59726 33406 59778 33458
rect 61406 33406 61458 33458
rect 62078 33406 62130 33458
rect 64206 33406 64258 33458
rect 68574 33406 68626 33458
rect 70478 33406 70530 33458
rect 72606 33406 72658 33458
rect 73502 33406 73554 33458
rect 81118 33406 81170 33458
rect 86494 33406 86546 33458
rect 88622 33406 88674 33458
rect 89518 33406 89570 33458
rect 91646 33406 91698 33458
rect 95342 33406 95394 33458
rect 97470 33406 97522 33458
rect 51662 33294 51714 33346
rect 54462 33294 54514 33346
rect 58382 33294 58434 33346
rect 59166 33294 59218 33346
rect 60398 33294 60450 33346
rect 64990 33294 65042 33346
rect 65774 33294 65826 33346
rect 69694 33294 69746 33346
rect 74286 33294 74338 33346
rect 74734 33294 74786 33346
rect 76302 33294 76354 33346
rect 78318 33294 78370 33346
rect 82798 33294 82850 33346
rect 83918 33294 83970 33346
rect 85822 33294 85874 33346
rect 92430 33294 92482 33346
rect 94558 33294 94610 33346
rect 51326 33182 51378 33234
rect 55246 33182 55298 33234
rect 58942 33182 58994 33234
rect 60622 33182 60674 33234
rect 66446 33182 66498 33234
rect 77310 33182 77362 33234
rect 77646 33182 77698 33234
rect 78990 33182 79042 33234
rect 82910 33182 82962 33234
rect 58046 33070 58098 33122
rect 73054 33070 73106 33122
rect 75742 33070 75794 33122
rect 81790 33070 81842 33122
rect 83582 33070 83634 33122
rect 84366 33070 84418 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 53790 32734 53842 32786
rect 54462 32734 54514 32786
rect 57822 32734 57874 32786
rect 58382 32734 58434 32786
rect 59726 32734 59778 32786
rect 60734 32734 60786 32786
rect 61070 32734 61122 32786
rect 61742 32734 61794 32786
rect 63534 32734 63586 32786
rect 71374 32734 71426 32786
rect 72606 32734 72658 32786
rect 73838 32734 73890 32786
rect 74286 32734 74338 32786
rect 75070 32734 75122 32786
rect 75518 32734 75570 32786
rect 76750 32734 76802 32786
rect 80670 32734 80722 32786
rect 81342 32734 81394 32786
rect 85598 32734 85650 32786
rect 86046 32734 86098 32786
rect 86718 32734 86770 32786
rect 88510 32734 88562 32786
rect 89182 32734 89234 32786
rect 94110 32734 94162 32786
rect 94670 32734 94722 32786
rect 95230 32734 95282 32786
rect 56590 32622 56642 32674
rect 62638 32622 62690 32674
rect 70254 32622 70306 32674
rect 76190 32622 76242 32674
rect 77870 32622 77922 32674
rect 81678 32622 81730 32674
rect 83022 32622 83074 32674
rect 87390 32622 87442 32674
rect 87838 32622 87890 32674
rect 90750 32622 90802 32674
rect 95790 32622 95842 32674
rect 96238 32622 96290 32674
rect 54798 32510 54850 32562
rect 55470 32510 55522 32562
rect 55806 32510 55858 32562
rect 56478 32510 56530 32562
rect 57598 32510 57650 32562
rect 62078 32510 62130 32562
rect 62862 32510 62914 32562
rect 65774 32510 65826 32562
rect 70366 32510 70418 32562
rect 70926 32510 70978 32562
rect 72046 32510 72098 32562
rect 73278 32510 73330 32562
rect 77086 32510 77138 32562
rect 77534 32510 77586 32562
rect 82350 32510 82402 32562
rect 90190 32510 90242 32562
rect 90974 32510 91026 32562
rect 91534 32510 91586 32562
rect 95566 32510 95618 32562
rect 66446 32398 66498 32450
rect 68574 32398 68626 32450
rect 69582 32398 69634 32450
rect 85150 32398 85202 32450
rect 69246 32286 69298 32338
rect 87054 32286 87106 32338
rect 89854 32286 89906 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 57038 31838 57090 31890
rect 57934 31838 57986 31890
rect 61406 31838 61458 31890
rect 68574 31838 68626 31890
rect 70366 31838 70418 31890
rect 71598 31838 71650 31890
rect 73726 31838 73778 31890
rect 76414 31838 76466 31890
rect 86942 31838 86994 31890
rect 89294 31838 89346 31890
rect 55918 31726 55970 31778
rect 67006 31726 67058 31778
rect 68014 31726 68066 31778
rect 70814 31726 70866 31778
rect 89854 31726 89906 31778
rect 55582 31614 55634 31666
rect 66670 31614 66722 31666
rect 67678 31614 67730 31666
rect 69358 31614 69410 31666
rect 69694 31614 69746 31666
rect 84142 31614 84194 31666
rect 90078 31614 90130 31666
rect 57374 31502 57426 31554
rect 83806 31502 83858 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 70590 31166 70642 31218
rect 83918 31054 83970 31106
rect 83134 30942 83186 30994
rect 69022 30830 69074 30882
rect 86046 30830 86098 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 83694 29598 83746 29650
rect 84254 29598 84306 29650
rect 85150 29486 85202 29538
rect 83246 29374 83298 29426
rect 84590 29374 84642 29426
rect 85374 29374 85426 29426
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 95230 25342 95282 25394
rect 94894 25230 94946 25282
rect 95790 25230 95842 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 1822 12798 1874 12850
rect 2158 12686 2210 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 1822 12350 1874 12402
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 6190 3390 6242 3442
rect 6638 3390 6690 3442
rect 18622 3390 18674 3442
rect 19070 3390 19122 3442
rect 31054 3390 31106 3442
rect 31502 3390 31554 3442
rect 44270 3390 44322 3442
rect 44942 3390 44994 3442
rect 56030 3390 56082 3442
rect 56702 3390 56754 3442
rect 67790 3390 67842 3442
rect 68798 3390 68850 3442
rect 80782 3390 80834 3442
rect 81230 3390 81282 3442
rect 93214 3390 93266 3442
rect 93998 3390 94050 3442
rect 6974 3278 7026 3330
rect 19406 3278 19458 3330
rect 31838 3278 31890 3330
rect 45278 3278 45330 3330
rect 57038 3278 57090 3330
rect 69134 3278 69186 3330
rect 81566 3278 81618 3330
rect 93662 3278 93714 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
<< metal2 >>
rect 6384 99200 6496 100000
rect 18816 99200 18928 100000
rect 31248 99200 31360 100000
rect 43680 99200 43792 100000
rect 56112 99200 56224 100000
rect 68544 99200 68656 100000
rect 80976 99200 81088 100000
rect 93408 99200 93520 100000
rect 6412 96628 6468 99200
rect 18844 97636 18900 99200
rect 18844 97580 19236 97636
rect 6412 96572 6804 96628
rect 4476 96460 4740 96470
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4476 96394 4740 96404
rect 6748 96178 6804 96572
rect 6748 96126 6750 96178
rect 6802 96126 6804 96178
rect 6748 96114 6804 96126
rect 19180 96178 19236 97580
rect 19180 96126 19182 96178
rect 19234 96126 19236 96178
rect 19180 96114 19236 96126
rect 31276 96178 31332 99200
rect 43708 96626 43764 99200
rect 43708 96574 43710 96626
rect 43762 96574 43764 96626
rect 43708 96562 43764 96574
rect 45052 96626 45108 96638
rect 45052 96574 45054 96626
rect 45106 96574 45108 96626
rect 35196 96460 35460 96470
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35196 96394 35460 96404
rect 31276 96126 31278 96178
rect 31330 96126 31332 96178
rect 31276 96114 31332 96126
rect 45052 96178 45108 96574
rect 56140 96626 56196 99200
rect 56140 96574 56142 96626
rect 56194 96574 56196 96626
rect 56140 96562 56196 96574
rect 56812 96626 56868 96638
rect 56812 96574 56814 96626
rect 56866 96574 56868 96626
rect 45052 96126 45054 96178
rect 45106 96126 45108 96178
rect 45052 96114 45108 96126
rect 56812 96178 56868 96574
rect 68572 96628 68628 99200
rect 81004 97636 81060 99200
rect 81004 97580 81396 97636
rect 68572 96572 68964 96628
rect 65916 96460 66180 96470
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 65916 96394 66180 96404
rect 56812 96126 56814 96178
rect 56866 96126 56868 96178
rect 56812 96114 56868 96126
rect 68908 96178 68964 96572
rect 68908 96126 68910 96178
rect 68962 96126 68964 96178
rect 68908 96114 68964 96126
rect 81340 96178 81396 97580
rect 81340 96126 81342 96178
rect 81394 96126 81396 96178
rect 81340 96114 81396 96126
rect 93436 96180 93492 99200
rect 96636 96460 96900 96470
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96636 96394 96900 96404
rect 93436 96114 93492 96124
rect 94332 96180 94388 96190
rect 94332 96086 94388 96124
rect 7868 96068 7924 96078
rect 7868 95974 7924 96012
rect 8316 96068 8372 96078
rect 8316 95974 8372 96012
rect 20300 96066 20356 96078
rect 20300 96014 20302 96066
rect 20354 96014 20356 96066
rect 20300 95844 20356 96014
rect 32172 96066 32228 96078
rect 32172 96014 32174 96066
rect 32226 96014 32228 96066
rect 20300 95778 20356 95788
rect 21308 95844 21364 95854
rect 21308 95750 21364 95788
rect 27692 95844 27748 95854
rect 19836 95676 20100 95686
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 19836 95610 20100 95620
rect 4476 94892 4740 94902
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4476 94826 4740 94836
rect 19836 94108 20100 94118
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 19836 94042 20100 94052
rect 4476 93324 4740 93334
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4476 93258 4740 93268
rect 19836 92540 20100 92550
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 19836 92474 20100 92484
rect 4476 91756 4740 91766
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4476 91690 4740 91700
rect 19836 90972 20100 90982
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 19836 90906 20100 90916
rect 4476 90188 4740 90198
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4476 90122 4740 90132
rect 19836 89404 20100 89414
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 19836 89338 20100 89348
rect 4476 88620 4740 88630
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4476 88554 4740 88564
rect 3276 88340 3332 88350
rect 3276 88246 3332 88284
rect 12572 88340 12628 88350
rect 1932 88116 1988 88126
rect 1708 88114 1988 88116
rect 1708 88062 1934 88114
rect 1986 88062 1988 88114
rect 1708 88060 1988 88062
rect 1708 87444 1764 88060
rect 1932 88050 1988 88060
rect 1708 87350 1764 87388
rect 4476 87052 4740 87062
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4476 86986 4740 86996
rect 4476 85484 4740 85494
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4476 85418 4740 85428
rect 4476 83916 4740 83926
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4476 83850 4740 83860
rect 4476 82348 4740 82358
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4476 82282 4740 82292
rect 4476 80780 4740 80790
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4476 80714 4740 80724
rect 4476 79212 4740 79222
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4476 79146 4740 79156
rect 4476 77644 4740 77654
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4476 77578 4740 77588
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 12572 63700 12628 88284
rect 19836 87836 20100 87846
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 19836 87770 20100 87780
rect 19836 86268 20100 86278
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 19836 86202 20100 86212
rect 19836 84700 20100 84710
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 19836 84634 20100 84644
rect 19836 83132 20100 83142
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 19836 83066 20100 83076
rect 19836 81564 20100 81574
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 19836 81498 20100 81508
rect 19836 79996 20100 80006
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 19836 79930 20100 79940
rect 19836 78428 20100 78438
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 19836 78362 20100 78372
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 27692 64820 27748 95788
rect 27692 64754 27748 64764
rect 32172 95844 32228 96014
rect 45948 96066 46004 96078
rect 45948 96014 45950 96066
rect 46002 96014 46004 96066
rect 33068 95844 33124 95854
rect 32172 95842 33124 95844
rect 32172 95790 33070 95842
rect 33122 95790 33124 95842
rect 32172 95788 33124 95790
rect 32172 64708 32228 95788
rect 33068 95778 33124 95788
rect 45948 95844 46004 96014
rect 47964 96068 48020 96078
rect 57708 96068 57764 96078
rect 58380 96068 58436 96078
rect 46620 95844 46676 95854
rect 45948 95842 46676 95844
rect 45948 95790 46622 95842
rect 46674 95790 46676 95842
rect 45948 95788 46676 95790
rect 35196 94892 35460 94902
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35196 94826 35460 94836
rect 35196 93324 35460 93334
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35196 93258 35460 93268
rect 35196 91756 35460 91766
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35196 91690 35460 91700
rect 35196 90188 35460 90198
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35196 90122 35460 90132
rect 35196 88620 35460 88630
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35196 88554 35460 88564
rect 35196 87052 35460 87062
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35196 86986 35460 86996
rect 35196 85484 35460 85494
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35196 85418 35460 85428
rect 35196 83916 35460 83926
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35196 83850 35460 83860
rect 35196 82348 35460 82358
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35196 82282 35460 82292
rect 35196 80780 35460 80790
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35196 80714 35460 80724
rect 35196 79212 35460 79222
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35196 79146 35460 79156
rect 35196 77644 35460 77654
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35196 77578 35460 77588
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 45948 68740 46004 95788
rect 46620 95778 46676 95788
rect 47852 70866 47908 70878
rect 47852 70814 47854 70866
rect 47906 70814 47908 70866
rect 47852 68964 47908 70814
rect 47852 68898 47908 68908
rect 45948 68674 46004 68684
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 32172 64642 32228 64652
rect 46956 64708 47012 64718
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 12572 63634 12628 63644
rect 46956 63588 47012 64652
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 46956 63522 47012 63532
rect 35196 63466 35460 63476
rect 47964 63252 48020 96012
rect 57596 96066 58436 96068
rect 57596 96014 57710 96066
rect 57762 96014 58382 96066
rect 58434 96014 58436 96066
rect 57596 96012 58436 96014
rect 50556 95676 50820 95686
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50556 95610 50820 95620
rect 50556 94108 50820 94118
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50556 94042 50820 94052
rect 50556 92540 50820 92550
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50556 92474 50820 92484
rect 50556 90972 50820 90982
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50556 90906 50820 90916
rect 50556 89404 50820 89414
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50556 89338 50820 89348
rect 54796 88002 54852 88014
rect 57372 88004 57428 88014
rect 54796 87950 54798 88002
rect 54850 87950 54852 88002
rect 50556 87836 50820 87846
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50556 87770 50820 87780
rect 54348 87554 54404 87566
rect 54348 87502 54350 87554
rect 54402 87502 54404 87554
rect 54236 87442 54292 87454
rect 54236 87390 54238 87442
rect 54290 87390 54292 87442
rect 54236 87332 54292 87390
rect 54236 87266 54292 87276
rect 53228 87220 53284 87230
rect 52556 87218 53284 87220
rect 52556 87166 53230 87218
rect 53282 87166 53284 87218
rect 52556 87164 53284 87166
rect 52556 86658 52612 87164
rect 53228 87154 53284 87164
rect 53564 87220 53620 87230
rect 53564 87126 53620 87164
rect 52556 86606 52558 86658
rect 52610 86606 52612 86658
rect 52556 86594 52612 86606
rect 53900 86660 53956 86670
rect 53900 86658 54068 86660
rect 53900 86606 53902 86658
rect 53954 86606 54068 86658
rect 53900 86604 54068 86606
rect 53900 86594 53956 86604
rect 52220 86436 52276 86446
rect 53564 86436 53620 86446
rect 51772 86434 52276 86436
rect 51772 86382 52222 86434
rect 52274 86382 52276 86434
rect 51772 86380 52276 86382
rect 50556 86268 50820 86278
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50556 86202 50820 86212
rect 51212 85874 51268 85886
rect 51212 85822 51214 85874
rect 51266 85822 51268 85874
rect 50556 84700 50820 84710
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50556 84634 50820 84644
rect 51100 84308 51156 84318
rect 51212 84308 51268 85822
rect 51772 84418 51828 86380
rect 52220 86370 52276 86380
rect 52556 86434 53620 86436
rect 52556 86382 53566 86434
rect 53618 86382 53620 86434
rect 52556 86380 53620 86382
rect 51884 85764 51940 85774
rect 51884 85762 52052 85764
rect 51884 85710 51886 85762
rect 51938 85710 52052 85762
rect 51884 85708 52052 85710
rect 51884 85698 51940 85708
rect 51996 85316 52052 85708
rect 51996 85260 52276 85316
rect 52220 84978 52276 85260
rect 52556 85090 52612 86380
rect 53564 86370 53620 86380
rect 54012 85988 54068 86604
rect 54012 85762 54068 85932
rect 54012 85710 54014 85762
rect 54066 85710 54068 85762
rect 54012 85698 54068 85710
rect 54348 86548 54404 87502
rect 54796 87332 54852 87950
rect 57148 88002 57428 88004
rect 57148 87950 57374 88002
rect 57426 87950 57428 88002
rect 57148 87948 57428 87950
rect 55580 87444 55636 87454
rect 55580 87442 55748 87444
rect 55580 87390 55582 87442
rect 55634 87390 55748 87442
rect 55580 87388 55748 87390
rect 55580 87378 55636 87388
rect 54796 87266 54852 87276
rect 55020 87332 55076 87342
rect 54684 86660 54740 86670
rect 55020 86660 55076 87276
rect 54684 86658 55076 86660
rect 54684 86606 54686 86658
rect 54738 86606 55076 86658
rect 54684 86604 55076 86606
rect 55580 86658 55636 86670
rect 55580 86606 55582 86658
rect 55634 86606 55636 86658
rect 54460 86548 54516 86558
rect 54348 86546 54516 86548
rect 54348 86494 54462 86546
rect 54514 86494 54516 86546
rect 54348 86492 54516 86494
rect 52556 85038 52558 85090
rect 52610 85038 52612 85090
rect 52556 85026 52612 85038
rect 52220 84926 52222 84978
rect 52274 84926 52276 84978
rect 52220 84914 52276 84926
rect 53788 84868 53844 84878
rect 53788 84774 53844 84812
rect 51772 84366 51774 84418
rect 51826 84366 51828 84418
rect 51772 84354 51828 84366
rect 51100 84306 51268 84308
rect 51100 84254 51102 84306
rect 51154 84254 51268 84306
rect 51100 84252 51268 84254
rect 51100 84242 51156 84252
rect 50556 83132 50820 83142
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50556 83066 50820 83076
rect 49756 81954 49812 81966
rect 49756 81902 49758 81954
rect 49810 81902 49812 81954
rect 49756 81172 49812 81902
rect 50540 81844 50596 81854
rect 50428 81842 50596 81844
rect 50428 81790 50542 81842
rect 50594 81790 50596 81842
rect 50428 81788 50596 81790
rect 50428 81396 50484 81788
rect 50540 81778 50596 81788
rect 50556 81564 50820 81574
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50556 81498 50820 81508
rect 50764 81396 50820 81406
rect 50428 81394 50820 81396
rect 50428 81342 50766 81394
rect 50818 81342 50820 81394
rect 50428 81340 50820 81342
rect 50764 81330 50820 81340
rect 50204 81284 50260 81294
rect 49532 80388 49588 80398
rect 49756 80388 49812 81116
rect 49532 80386 49812 80388
rect 49532 80334 49534 80386
rect 49586 80334 49812 80386
rect 49532 80332 49812 80334
rect 49980 81282 50260 81284
rect 49980 81230 50206 81282
rect 50258 81230 50260 81282
rect 49980 81228 50260 81230
rect 49532 79602 49588 80332
rect 49532 79550 49534 79602
rect 49586 79550 49588 79602
rect 49532 79538 49588 79550
rect 49308 78708 49364 78718
rect 49308 78614 49364 78652
rect 49756 78596 49812 78606
rect 49644 78540 49756 78596
rect 48860 78260 48916 78270
rect 48860 78166 48916 78204
rect 49644 78260 49700 78540
rect 49756 78502 49812 78540
rect 48300 78148 48356 78158
rect 48300 78054 48356 78092
rect 49644 78146 49700 78204
rect 49980 78258 50036 81228
rect 50204 81218 50260 81228
rect 50316 81284 50372 81294
rect 50988 81284 51044 81294
rect 50316 81190 50372 81228
rect 50876 81282 51044 81284
rect 50876 81230 50990 81282
rect 51042 81230 51044 81282
rect 50876 81228 51044 81230
rect 50204 80948 50260 80958
rect 50204 80946 50372 80948
rect 50204 80894 50206 80946
rect 50258 80894 50372 80946
rect 50204 80892 50372 80894
rect 50204 80882 50260 80892
rect 50204 80274 50260 80286
rect 50204 80222 50206 80274
rect 50258 80222 50260 80274
rect 50204 78820 50260 80222
rect 50316 79714 50372 80892
rect 50556 79996 50820 80006
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50556 79930 50820 79940
rect 50316 79662 50318 79714
rect 50370 79662 50372 79714
rect 50316 79650 50372 79662
rect 50204 78754 50260 78764
rect 49980 78206 49982 78258
rect 50034 78206 50036 78258
rect 49980 78194 50036 78206
rect 50092 78708 50148 78718
rect 49644 78094 49646 78146
rect 49698 78094 49700 78146
rect 49644 78082 49700 78094
rect 49756 78148 49812 78158
rect 49756 78054 49812 78092
rect 50092 77364 50148 78652
rect 50652 78706 50708 78718
rect 50652 78654 50654 78706
rect 50706 78654 50708 78706
rect 50204 78596 50260 78606
rect 50652 78596 50708 78654
rect 50764 78708 50820 78718
rect 50764 78614 50820 78652
rect 50260 78540 50708 78596
rect 50204 78464 50260 78540
rect 50428 78260 50484 78540
rect 50556 78428 50820 78438
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50556 78362 50820 78372
rect 50092 77298 50148 77308
rect 50316 78148 50372 78158
rect 49868 77250 49924 77262
rect 49868 77198 49870 77250
rect 49922 77198 49924 77250
rect 49868 77028 49924 77198
rect 49868 75682 49924 76972
rect 49868 75630 49870 75682
rect 49922 75630 49924 75682
rect 49868 74900 49924 75630
rect 50316 75572 50372 78092
rect 50428 78146 50484 78204
rect 50764 78260 50820 78270
rect 50876 78260 50932 81228
rect 50988 81218 51044 81228
rect 51100 81170 51156 81182
rect 51100 81118 51102 81170
rect 51154 81118 51156 81170
rect 51100 80948 51156 81118
rect 51212 81172 51268 84252
rect 53900 84196 53956 84206
rect 54348 84196 54404 86492
rect 54460 86482 54516 86492
rect 54684 86100 54740 86604
rect 55356 86436 55412 86446
rect 54684 86034 54740 86044
rect 55132 86434 55412 86436
rect 55132 86382 55358 86434
rect 55410 86382 55412 86434
rect 55132 86380 55412 86382
rect 54572 85762 54628 85774
rect 54572 85710 54574 85762
rect 54626 85710 54628 85762
rect 54460 85090 54516 85102
rect 54460 85038 54462 85090
rect 54514 85038 54516 85090
rect 54460 84868 54516 85038
rect 54460 84756 54516 84812
rect 54572 84756 54628 85710
rect 55132 85202 55188 86380
rect 55356 86370 55412 86380
rect 55468 86100 55524 86110
rect 55580 86100 55636 86606
rect 55468 86098 55636 86100
rect 55468 86046 55470 86098
rect 55522 86046 55636 86098
rect 55468 86044 55636 86046
rect 55468 86034 55524 86044
rect 55692 85988 55748 87388
rect 56028 87442 56084 87454
rect 56028 87390 56030 87442
rect 56082 87390 56084 87442
rect 56028 87220 56084 87390
rect 56028 87154 56084 87164
rect 56476 86772 56532 86782
rect 56476 86658 56532 86716
rect 57148 86770 57204 87948
rect 57372 87938 57428 87948
rect 57484 87330 57540 87342
rect 57484 87278 57486 87330
rect 57538 87278 57540 87330
rect 57484 87220 57540 87278
rect 57484 87154 57540 87164
rect 57596 86996 57652 96012
rect 57708 96002 57764 96012
rect 58380 96002 58436 96012
rect 70028 96066 70084 96078
rect 70028 96014 70030 96066
rect 70082 96014 70084 96066
rect 70028 95844 70084 96014
rect 82348 96066 82404 96078
rect 82348 96014 82350 96066
rect 82402 96014 82404 96066
rect 70028 95778 70084 95788
rect 70476 95844 70532 95854
rect 70476 95750 70532 95788
rect 77980 95844 78036 95854
rect 65916 94892 66180 94902
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 65916 94826 66180 94836
rect 65916 93324 66180 93334
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 65916 93258 66180 93268
rect 65916 91756 66180 91766
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 65916 91690 66180 91700
rect 77980 90748 78036 95788
rect 82348 95844 82404 96014
rect 93100 96068 93156 96078
rect 93100 95974 93156 96012
rect 93884 96068 93940 96078
rect 93884 95974 93940 96012
rect 97468 96068 97524 96078
rect 82908 95844 82964 95854
rect 82348 95842 82964 95844
rect 82348 95790 82910 95842
rect 82962 95790 82964 95842
rect 82348 95788 82964 95790
rect 81276 95676 81540 95686
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81276 95610 81540 95620
rect 81276 94108 81540 94118
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81276 94042 81540 94052
rect 81276 92540 81540 92550
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81276 92474 81540 92484
rect 81276 90972 81540 90982
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81276 90906 81540 90916
rect 77980 90692 78484 90748
rect 65916 90188 66180 90198
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 65916 90122 66180 90132
rect 68236 89010 68292 89022
rect 68236 88958 68238 89010
rect 68290 88958 68292 89010
rect 63084 88898 63140 88910
rect 63532 88900 63588 88910
rect 63084 88846 63086 88898
rect 63138 88846 63140 88898
rect 61852 88226 61908 88238
rect 61852 88174 61854 88226
rect 61906 88174 61908 88226
rect 57708 88114 57764 88126
rect 57708 88062 57710 88114
rect 57762 88062 57764 88114
rect 57708 87668 57764 88062
rect 59612 88002 59668 88014
rect 60620 88004 60676 88014
rect 59612 87950 59614 88002
rect 59666 87950 59668 88002
rect 59052 87892 59108 87902
rect 58044 87668 58100 87678
rect 57708 87666 58100 87668
rect 57708 87614 58046 87666
rect 58098 87614 58100 87666
rect 57708 87612 58100 87614
rect 58044 87602 58100 87612
rect 59052 87442 59108 87836
rect 59612 87892 59668 87950
rect 60508 88002 60676 88004
rect 60508 87950 60622 88002
rect 60674 87950 60676 88002
rect 60508 87948 60676 87950
rect 59612 87826 59668 87836
rect 60284 87892 60340 87902
rect 59164 87556 59220 87566
rect 59164 87554 59332 87556
rect 59164 87502 59166 87554
rect 59218 87502 59332 87554
rect 59164 87500 59332 87502
rect 59164 87490 59220 87500
rect 59052 87390 59054 87442
rect 59106 87390 59108 87442
rect 57596 86930 57652 86940
rect 57820 87220 57876 87230
rect 57148 86718 57150 86770
rect 57202 86718 57204 86770
rect 57148 86706 57204 86718
rect 57596 86772 57652 86782
rect 56476 86606 56478 86658
rect 56530 86606 56532 86658
rect 56476 86594 56532 86606
rect 55692 85922 55748 85932
rect 56476 86100 56532 86110
rect 56476 85874 56532 86044
rect 56476 85822 56478 85874
rect 56530 85822 56532 85874
rect 56476 85810 56532 85822
rect 56588 85986 56644 85998
rect 56588 85934 56590 85986
rect 56642 85934 56644 85986
rect 55132 85150 55134 85202
rect 55186 85150 55188 85202
rect 55132 85138 55188 85150
rect 55804 85764 55860 85774
rect 54460 84700 54628 84756
rect 53900 84194 54404 84196
rect 53900 84142 53902 84194
rect 53954 84142 54404 84194
rect 53900 84140 54404 84142
rect 54460 84194 54516 84206
rect 54460 84142 54462 84194
rect 54514 84142 54516 84194
rect 53900 84130 53956 84140
rect 53228 83636 53284 83646
rect 52444 83300 52500 83310
rect 52220 82740 52276 82750
rect 51212 81106 51268 81116
rect 51660 81172 51716 81182
rect 51660 81078 51716 81116
rect 51100 80882 51156 80892
rect 52108 78820 52164 78830
rect 52108 78726 52164 78764
rect 51660 78706 51716 78718
rect 51660 78654 51662 78706
rect 51714 78654 51716 78706
rect 50988 78596 51044 78606
rect 51324 78596 51380 78606
rect 51548 78596 51604 78606
rect 50988 78502 51044 78540
rect 51100 78594 51380 78596
rect 51100 78542 51326 78594
rect 51378 78542 51380 78594
rect 51100 78540 51380 78542
rect 50764 78258 50932 78260
rect 50764 78206 50766 78258
rect 50818 78206 50932 78258
rect 50764 78204 50932 78206
rect 50764 78194 50820 78204
rect 50428 78094 50430 78146
rect 50482 78094 50484 78146
rect 50428 78082 50484 78094
rect 50540 78146 50596 78158
rect 50540 78094 50542 78146
rect 50594 78094 50596 78146
rect 50540 78036 50596 78094
rect 50540 77970 50596 77980
rect 51100 77364 51156 78540
rect 51324 78530 51380 78540
rect 51436 78594 51604 78596
rect 51436 78542 51550 78594
rect 51602 78542 51604 78594
rect 51436 78540 51604 78542
rect 51324 78148 51380 78158
rect 51324 78054 51380 78092
rect 51212 78034 51268 78046
rect 51212 77982 51214 78034
rect 51266 77982 51268 78034
rect 51212 77924 51268 77982
rect 51212 77858 51268 77868
rect 50428 77308 51156 77364
rect 50428 75796 50484 77308
rect 50540 77140 50596 77150
rect 50540 77138 51380 77140
rect 50540 77086 50542 77138
rect 50594 77086 51380 77138
rect 50540 77084 51380 77086
rect 50540 77074 50596 77084
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50876 76356 50932 76366
rect 50652 76354 50932 76356
rect 50652 76302 50878 76354
rect 50930 76302 50932 76354
rect 50652 76300 50932 76302
rect 50540 75796 50596 75806
rect 50428 75794 50596 75796
rect 50428 75742 50542 75794
rect 50594 75742 50596 75794
rect 50428 75740 50596 75742
rect 50540 75730 50596 75740
rect 50652 75572 50708 76300
rect 50876 76290 50932 76300
rect 50316 75516 50708 75572
rect 49980 74900 50036 74910
rect 49868 74898 50036 74900
rect 49868 74846 49982 74898
rect 50034 74846 50036 74898
rect 49868 74844 50036 74846
rect 49980 74834 50036 74844
rect 50204 74228 50260 74238
rect 50204 74134 50260 74172
rect 49756 72546 49812 72558
rect 49756 72494 49758 72546
rect 49810 72494 49812 72546
rect 49756 71988 49812 72494
rect 49756 71922 49812 71932
rect 49980 72322 50036 72334
rect 49980 72270 49982 72322
rect 50034 72270 50036 72322
rect 48860 70980 48916 70990
rect 48860 70978 49028 70980
rect 48860 70926 48862 70978
rect 48914 70926 49028 70978
rect 48860 70924 49028 70926
rect 48860 70914 48916 70924
rect 48188 70868 48244 70878
rect 48188 70774 48244 70812
rect 47964 63186 48020 63196
rect 48076 70756 48132 70766
rect 1820 63026 1876 63038
rect 1820 62974 1822 63026
rect 1874 62974 1876 63026
rect 1820 62468 1876 62974
rect 2156 62914 2212 62926
rect 2156 62862 2158 62914
rect 2210 62862 2212 62914
rect 2156 62804 2212 62862
rect 2156 62738 2212 62748
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 1820 62374 1876 62412
rect 47852 62242 47908 62254
rect 47852 62190 47854 62242
rect 47906 62190 47908 62242
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 47852 61796 47908 62190
rect 48076 61796 48132 70700
rect 48972 69412 49028 70924
rect 49532 70868 49588 70878
rect 49532 70774 49588 70812
rect 48972 67842 49028 69356
rect 49532 69412 49588 69422
rect 49532 69318 49588 69356
rect 49980 69300 50036 72270
rect 50316 69636 50372 75516
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50764 75012 50820 75022
rect 50764 74918 50820 74956
rect 50652 74228 50708 74238
rect 50652 74114 50708 74172
rect 50652 74062 50654 74114
rect 50706 74062 50708 74114
rect 50652 74050 50708 74062
rect 51324 74114 51380 77084
rect 51324 74062 51326 74114
rect 51378 74062 51380 74114
rect 51324 74050 51380 74062
rect 50988 74004 51044 74014
rect 50988 74002 51268 74004
rect 50988 73950 50990 74002
rect 51042 73950 51268 74002
rect 50988 73948 51268 73950
rect 51436 73948 51492 78540
rect 51548 78530 51604 78540
rect 50988 73938 51044 73948
rect 50764 73892 50820 73902
rect 51212 73892 51492 73948
rect 51548 78034 51604 78046
rect 51548 77982 51550 78034
rect 51602 77982 51604 78034
rect 50764 73890 50932 73892
rect 50764 73838 50766 73890
rect 50818 73838 50932 73890
rect 50764 73836 50932 73838
rect 50764 73826 50820 73836
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50876 73220 50932 73836
rect 51548 73890 51604 77982
rect 51660 77140 51716 78654
rect 52220 78260 52276 82684
rect 52444 81282 52500 83244
rect 52668 83300 52724 83310
rect 52668 83298 52836 83300
rect 52668 83246 52670 83298
rect 52722 83246 52836 83298
rect 52668 83244 52836 83246
rect 52668 83234 52724 83244
rect 52668 82068 52724 82078
rect 52668 81974 52724 82012
rect 52780 81956 52836 83244
rect 52892 82740 52948 82750
rect 52892 82646 52948 82684
rect 52780 81890 52836 81900
rect 52444 81230 52446 81282
rect 52498 81230 52500 81282
rect 52444 81218 52500 81230
rect 52332 80500 52388 80510
rect 52332 80498 53172 80500
rect 52332 80446 52334 80498
rect 52386 80446 53172 80498
rect 52332 80444 53172 80446
rect 52332 80434 52388 80444
rect 52332 79828 52388 79838
rect 52332 78988 52388 79772
rect 52892 79828 52948 79838
rect 52892 79734 52948 79772
rect 53116 79826 53172 80444
rect 53116 79774 53118 79826
rect 53170 79774 53172 79826
rect 53116 79762 53172 79774
rect 53228 80164 53284 83580
rect 53676 83636 53732 83646
rect 53676 83522 53732 83580
rect 54460 83636 54516 84142
rect 54572 84196 54628 84700
rect 54796 84196 54852 84206
rect 55804 84196 55860 85708
rect 56588 85204 56644 85934
rect 56588 85138 56644 85148
rect 56700 85988 56756 85998
rect 54572 84194 54964 84196
rect 54572 84142 54798 84194
rect 54850 84142 54964 84194
rect 54572 84140 54964 84142
rect 54796 84130 54852 84140
rect 54460 83570 54516 83580
rect 53676 83470 53678 83522
rect 53730 83470 53732 83522
rect 53676 83458 53732 83470
rect 54460 83410 54516 83422
rect 54460 83358 54462 83410
rect 54514 83358 54516 83410
rect 53340 83300 53396 83310
rect 53340 83298 53508 83300
rect 53340 83246 53342 83298
rect 53394 83246 53508 83298
rect 53340 83244 53508 83246
rect 53340 83234 53396 83244
rect 53340 81956 53396 81966
rect 53340 81730 53396 81900
rect 53340 81678 53342 81730
rect 53394 81678 53396 81730
rect 53340 81172 53396 81678
rect 53340 80388 53396 81116
rect 53452 80948 53508 83244
rect 53564 83298 53620 83310
rect 53564 83246 53566 83298
rect 53618 83246 53620 83298
rect 53564 82068 53620 83246
rect 54124 83300 54180 83310
rect 54124 83206 54180 83244
rect 54348 83298 54404 83310
rect 54348 83246 54350 83298
rect 54402 83246 54404 83298
rect 53564 82002 53620 82012
rect 54124 82626 54180 82638
rect 54124 82574 54126 82626
rect 54178 82574 54180 82626
rect 54124 82292 54180 82574
rect 54124 81956 54180 82236
rect 54124 81862 54180 81900
rect 53452 80882 53508 80892
rect 54012 81284 54068 81294
rect 54012 80836 54068 81228
rect 54348 80836 54404 83246
rect 54012 80780 54404 80836
rect 53452 80388 53508 80398
rect 53340 80386 53732 80388
rect 53340 80334 53454 80386
rect 53506 80334 53732 80386
rect 53340 80332 53732 80334
rect 53452 80322 53508 80332
rect 53228 79714 53284 80108
rect 53676 79828 53732 80332
rect 54012 79940 54068 80780
rect 54460 80724 54516 83358
rect 54908 83298 54964 84140
rect 55804 84130 55860 84140
rect 56476 84196 56532 84206
rect 54908 83246 54910 83298
rect 54962 83246 54964 83298
rect 54908 82292 54964 83246
rect 54964 82236 55076 82292
rect 54908 82226 54964 82236
rect 54908 81842 54964 81854
rect 54908 81790 54910 81842
rect 54962 81790 54964 81842
rect 54908 81396 54964 81790
rect 55020 81732 55076 82236
rect 55020 81666 55076 81676
rect 54908 81340 55188 81396
rect 55020 81172 55076 81182
rect 54908 81170 55076 81172
rect 54908 81118 55022 81170
rect 55074 81118 55076 81170
rect 54908 81116 55076 81118
rect 54124 80668 54516 80724
rect 54572 81058 54628 81070
rect 54572 81006 54574 81058
rect 54626 81006 54628 81058
rect 54124 80276 54180 80668
rect 54236 80500 54292 80510
rect 54236 80406 54292 80444
rect 54124 80220 54404 80276
rect 54012 79884 54292 79940
rect 53676 79826 54180 79828
rect 53676 79774 53678 79826
rect 53730 79774 54180 79826
rect 53676 79772 54180 79774
rect 53676 79762 53732 79772
rect 53228 79662 53230 79714
rect 53282 79662 53284 79714
rect 52444 79492 52500 79502
rect 52444 79490 52612 79492
rect 52444 79438 52446 79490
rect 52498 79438 52612 79490
rect 52444 79436 52612 79438
rect 52444 79426 52500 79436
rect 52556 78988 52612 79436
rect 53228 79156 53284 79662
rect 53228 79100 53732 79156
rect 53676 79044 53732 79100
rect 52332 78932 52500 78988
rect 52556 78932 53620 78988
rect 52444 78818 52500 78932
rect 52444 78766 52446 78818
rect 52498 78766 52500 78818
rect 52444 78754 52500 78766
rect 53340 78820 53396 78830
rect 53340 78726 53396 78764
rect 53564 78706 53620 78932
rect 53564 78654 53566 78706
rect 53618 78654 53620 78706
rect 53564 78642 53620 78654
rect 53676 78706 53732 78988
rect 53676 78654 53678 78706
rect 53730 78654 53732 78706
rect 52332 78596 52388 78606
rect 52332 78502 52388 78540
rect 52220 78204 52388 78260
rect 52108 78146 52164 78158
rect 52108 78094 52110 78146
rect 52162 78094 52164 78146
rect 51660 77074 51716 77084
rect 51772 78036 51828 78046
rect 51660 75236 51716 75246
rect 51660 74114 51716 75180
rect 51660 74062 51662 74114
rect 51714 74062 51716 74114
rect 51660 74050 51716 74062
rect 51548 73838 51550 73890
rect 51602 73838 51604 73890
rect 51548 73826 51604 73838
rect 51324 73220 51380 73230
rect 51772 73220 51828 77980
rect 51884 78034 51940 78046
rect 52108 78036 52164 78094
rect 51884 77982 51886 78034
rect 51938 77982 51940 78034
rect 51884 75012 51940 77982
rect 51996 77980 52164 78036
rect 52220 78034 52276 78046
rect 52220 77982 52222 78034
rect 52274 77982 52276 78034
rect 51996 77588 52052 77980
rect 51996 77532 52164 77588
rect 51884 74946 51940 74956
rect 51996 77364 52052 77374
rect 51996 73948 52052 77308
rect 52108 74114 52164 77532
rect 52220 75124 52276 77982
rect 52332 77252 52388 78204
rect 53676 78258 53732 78654
rect 53676 78206 53678 78258
rect 53730 78206 53732 78258
rect 53676 78194 53732 78206
rect 54124 78258 54180 79772
rect 54236 78820 54292 79884
rect 54348 79826 54404 80220
rect 54348 79774 54350 79826
rect 54402 79774 54404 79826
rect 54348 79762 54404 79774
rect 54572 79716 54628 81006
rect 54908 80500 54964 81116
rect 55020 81106 55076 81116
rect 54908 80434 54964 80444
rect 55020 80948 55076 80958
rect 54572 79622 54628 79660
rect 54684 79604 54740 79614
rect 55020 79604 55076 80892
rect 55132 79826 55188 81340
rect 55132 79774 55134 79826
rect 55186 79774 55188 79826
rect 55132 79762 55188 79774
rect 55244 81282 55300 81294
rect 55244 81230 55246 81282
rect 55298 81230 55300 81282
rect 55244 79828 55300 81230
rect 56028 81282 56084 81294
rect 56028 81230 56030 81282
rect 56082 81230 56084 81282
rect 55356 81170 55412 81182
rect 55804 81172 55860 81182
rect 55356 81118 55358 81170
rect 55410 81118 55412 81170
rect 55356 80388 55412 81118
rect 55356 80322 55412 80332
rect 55468 81170 55860 81172
rect 55468 81118 55806 81170
rect 55858 81118 55860 81170
rect 55468 81116 55860 81118
rect 55244 79762 55300 79772
rect 55356 79714 55412 79726
rect 55356 79662 55358 79714
rect 55410 79662 55412 79714
rect 55356 79604 55412 79662
rect 55468 79714 55524 81116
rect 55804 81106 55860 81116
rect 56028 80612 56084 81230
rect 56028 80546 56084 80556
rect 56140 81170 56196 81182
rect 56140 81118 56142 81170
rect 56194 81118 56196 81170
rect 56140 80276 56196 81118
rect 56364 80500 56420 80510
rect 56364 80406 56420 80444
rect 55468 79662 55470 79714
rect 55522 79662 55524 79714
rect 55468 79650 55524 79662
rect 55916 80220 56140 80276
rect 55916 79826 55972 80220
rect 56140 80210 56196 80220
rect 55916 79774 55918 79826
rect 55970 79774 55972 79826
rect 55020 79548 55412 79604
rect 55916 79604 55972 79774
rect 54684 79510 54740 79548
rect 55916 79538 55972 79548
rect 54572 79044 54628 79054
rect 54572 78930 54628 78988
rect 54572 78878 54574 78930
rect 54626 78878 54628 78930
rect 54572 78866 54628 78878
rect 54236 78754 54292 78764
rect 54124 78206 54126 78258
rect 54178 78206 54180 78258
rect 54124 78194 54180 78206
rect 54236 78594 54292 78606
rect 54236 78542 54238 78594
rect 54290 78542 54292 78594
rect 52668 78036 52724 78046
rect 52668 77942 52724 77980
rect 53116 77924 53172 77934
rect 52332 77186 52388 77196
rect 52668 77362 52724 77374
rect 52668 77310 52670 77362
rect 52722 77310 52724 77362
rect 52668 76244 52724 77310
rect 52892 77252 52948 77262
rect 52892 76466 52948 77196
rect 52892 76414 52894 76466
rect 52946 76414 52948 76466
rect 52892 76402 52948 76414
rect 52668 76178 52724 76188
rect 52668 75794 52724 75806
rect 52668 75742 52670 75794
rect 52722 75742 52724 75794
rect 52668 75460 52724 75742
rect 52668 75394 52724 75404
rect 52220 75058 52276 75068
rect 52892 75012 52948 75022
rect 52892 74786 52948 74956
rect 52892 74734 52894 74786
rect 52946 74734 52948 74786
rect 52892 74722 52948 74734
rect 52108 74062 52110 74114
rect 52162 74062 52164 74114
rect 52108 74050 52164 74062
rect 52444 74228 52500 74238
rect 52444 74114 52500 74172
rect 53116 74228 53172 77868
rect 54236 77140 54292 78542
rect 54908 78148 54964 78158
rect 54796 78146 54964 78148
rect 54796 78094 54910 78146
rect 54962 78094 54964 78146
rect 54796 78092 54964 78094
rect 53340 77028 53396 77038
rect 53340 76934 53396 76972
rect 53788 77028 53844 77038
rect 53788 76356 53844 76972
rect 54236 76580 54292 77084
rect 54348 77250 54404 77262
rect 54348 77198 54350 77250
rect 54402 77198 54404 77250
rect 54348 77028 54404 77198
rect 54348 76962 54404 76972
rect 54236 76514 54292 76524
rect 53564 76244 53620 76254
rect 53340 75236 53396 75246
rect 53340 75122 53396 75180
rect 53340 75070 53342 75122
rect 53394 75070 53396 75122
rect 53340 75058 53396 75070
rect 53564 75122 53620 76188
rect 53788 75684 53844 76300
rect 53788 75682 53956 75684
rect 53788 75630 53790 75682
rect 53842 75630 53956 75682
rect 53788 75628 53956 75630
rect 53788 75618 53844 75628
rect 53564 75070 53566 75122
rect 53618 75070 53620 75122
rect 53564 75058 53620 75070
rect 53676 74898 53732 74910
rect 53676 74846 53678 74898
rect 53730 74846 53732 74898
rect 53676 74788 53732 74846
rect 53676 74722 53732 74732
rect 53116 74162 53172 74172
rect 53340 74228 53396 74238
rect 53340 74134 53396 74172
rect 53900 74226 53956 75628
rect 54572 75570 54628 75582
rect 54572 75518 54574 75570
rect 54626 75518 54628 75570
rect 54124 75124 54180 75134
rect 54124 74900 54180 75068
rect 54572 75124 54628 75518
rect 54796 75236 54852 78092
rect 54908 78082 54964 78092
rect 55020 78036 55076 78046
rect 56364 78036 56420 78046
rect 55020 78034 55300 78036
rect 55020 77982 55022 78034
rect 55074 77982 55300 78034
rect 55020 77980 55300 77982
rect 55020 77970 55076 77980
rect 54908 77812 54964 77822
rect 54908 77810 55188 77812
rect 54908 77758 54910 77810
rect 54962 77758 55188 77810
rect 54908 77756 55188 77758
rect 54908 77746 54964 77756
rect 55132 77362 55188 77756
rect 55132 77310 55134 77362
rect 55186 77310 55188 77362
rect 55132 77298 55188 77310
rect 55244 76692 55300 77980
rect 55244 76626 55300 76636
rect 56028 78034 56420 78036
rect 56028 77982 56366 78034
rect 56418 77982 56420 78034
rect 56028 77980 56420 77982
rect 54796 75170 54852 75180
rect 54908 76580 54964 76590
rect 54572 75058 54628 75068
rect 54908 75122 54964 76524
rect 54908 75070 54910 75122
rect 54962 75070 54964 75122
rect 54908 75058 54964 75070
rect 55132 75460 55188 75470
rect 55132 75122 55188 75404
rect 55132 75070 55134 75122
rect 55186 75070 55188 75122
rect 55132 75058 55188 75070
rect 55692 75124 55748 75134
rect 55692 75030 55748 75068
rect 54348 75012 54404 75022
rect 54348 74918 54404 74956
rect 55916 75010 55972 75022
rect 55916 74958 55918 75010
rect 55970 74958 55972 75010
rect 54124 74834 54180 74844
rect 54460 74898 54516 74910
rect 54460 74846 54462 74898
rect 54514 74846 54516 74898
rect 54460 74788 54516 74846
rect 55244 74898 55300 74910
rect 55244 74846 55246 74898
rect 55298 74846 55300 74898
rect 53900 74174 53902 74226
rect 53954 74174 53956 74226
rect 53900 74162 53956 74174
rect 54348 74228 54404 74238
rect 54460 74228 54516 74732
rect 54348 74226 54516 74228
rect 54348 74174 54350 74226
rect 54402 74174 54516 74226
rect 54348 74172 54516 74174
rect 54796 74788 54852 74798
rect 54796 74226 54852 74732
rect 55244 74788 55300 74846
rect 55916 74900 55972 74958
rect 56028 75010 56084 77980
rect 56364 77970 56420 77980
rect 56476 76580 56532 84140
rect 56588 81732 56644 81742
rect 56588 81394 56644 81676
rect 56588 81342 56590 81394
rect 56642 81342 56644 81394
rect 56588 81330 56644 81342
rect 56700 79828 56756 85932
rect 57596 85874 57652 86716
rect 57596 85822 57598 85874
rect 57650 85822 57652 85874
rect 57260 85204 57316 85214
rect 57260 85110 57316 85148
rect 56924 84308 56980 84318
rect 56924 83298 56980 84252
rect 57372 84196 57428 84206
rect 57372 84102 57428 84140
rect 56924 83246 56926 83298
rect 56978 83246 56980 83298
rect 56924 82740 56980 83246
rect 56924 82674 56980 82684
rect 57596 82738 57652 85822
rect 57708 86100 57764 86110
rect 57708 85202 57764 86044
rect 57708 85150 57710 85202
rect 57762 85150 57764 85202
rect 57708 85138 57764 85150
rect 57596 82686 57598 82738
rect 57650 82686 57652 82738
rect 57596 82674 57652 82686
rect 57036 82068 57092 82078
rect 56924 82066 57092 82068
rect 56924 82014 57038 82066
rect 57090 82014 57092 82066
rect 56924 82012 57092 82014
rect 56924 80612 56980 82012
rect 57036 82002 57092 82012
rect 56812 80388 56868 80398
rect 56812 80294 56868 80332
rect 56700 79734 56756 79772
rect 56028 74958 56030 75010
rect 56082 74958 56084 75010
rect 56028 74946 56084 74958
rect 56364 76524 56532 76580
rect 56588 79604 56644 79614
rect 56588 78146 56644 79548
rect 56924 79380 56980 80556
rect 57372 81058 57428 81070
rect 57372 81006 57374 81058
rect 57426 81006 57428 81058
rect 57036 80500 57092 80510
rect 57036 80274 57092 80444
rect 57148 80388 57204 80398
rect 57148 80294 57204 80332
rect 57372 80388 57428 81006
rect 57372 80322 57428 80332
rect 57484 80500 57540 80510
rect 57036 80222 57038 80274
rect 57090 80222 57092 80274
rect 57036 80210 57092 80222
rect 56924 79314 56980 79324
rect 57372 79716 57428 79726
rect 57372 78930 57428 79660
rect 57484 79714 57540 80444
rect 57596 80388 57652 80398
rect 57596 80294 57652 80332
rect 57484 79662 57486 79714
rect 57538 79662 57540 79714
rect 57484 79650 57540 79662
rect 57820 78988 57876 87164
rect 58380 87220 58436 87230
rect 58380 87126 58436 87164
rect 58716 86324 58772 86334
rect 58268 85988 58324 85998
rect 58268 85894 58324 85932
rect 58716 84978 58772 86268
rect 58716 84926 58718 84978
rect 58770 84926 58772 84978
rect 58716 84914 58772 84926
rect 59052 84978 59108 87390
rect 59276 86770 59332 87500
rect 59276 86718 59278 86770
rect 59330 86718 59332 86770
rect 59276 86324 59332 86718
rect 59948 87442 60004 87454
rect 59948 87390 59950 87442
rect 60002 87390 60004 87442
rect 59948 86772 60004 87390
rect 59948 86706 60004 86716
rect 60060 86658 60116 86670
rect 60060 86606 60062 86658
rect 60114 86606 60116 86658
rect 59276 86258 59332 86268
rect 59836 86434 59892 86446
rect 59836 86382 59838 86434
rect 59890 86382 59892 86434
rect 59836 85988 59892 86382
rect 59836 85922 59892 85932
rect 60060 85764 60116 86606
rect 59724 85708 60116 85764
rect 59388 85316 59444 85326
rect 59388 85222 59444 85260
rect 59724 85314 59780 85708
rect 59724 85262 59726 85314
rect 59778 85262 59780 85314
rect 59724 85250 59780 85262
rect 59052 84926 59054 84978
rect 59106 84926 59108 84978
rect 59052 84914 59108 84926
rect 59500 85204 59556 85214
rect 58828 84308 58884 84318
rect 58828 84214 58884 84252
rect 57932 83524 57988 83534
rect 57932 83522 58660 83524
rect 57932 83470 57934 83522
rect 57986 83470 58660 83522
rect 57932 83468 58660 83470
rect 57932 83458 57988 83468
rect 58156 83298 58212 83310
rect 58156 83246 58158 83298
rect 58210 83246 58212 83298
rect 58156 82852 58212 83246
rect 58268 82852 58324 82862
rect 58156 82850 58324 82852
rect 58156 82798 58270 82850
rect 58322 82798 58324 82850
rect 58156 82796 58324 82798
rect 58268 82786 58324 82796
rect 58604 82178 58660 83468
rect 58604 82126 58606 82178
rect 58658 82126 58660 82178
rect 58604 82114 58660 82126
rect 58940 82628 58996 82638
rect 58940 81954 58996 82572
rect 58940 81902 58942 81954
rect 58994 81902 58996 81954
rect 58492 79714 58548 79726
rect 58492 79662 58494 79714
rect 58546 79662 58548 79714
rect 57932 79602 57988 79614
rect 57932 79550 57934 79602
rect 57986 79550 57988 79602
rect 57932 79492 57988 79550
rect 58268 79604 58324 79614
rect 58268 79510 58324 79548
rect 57932 79426 57988 79436
rect 57820 78932 57988 78988
rect 57372 78878 57374 78930
rect 57426 78878 57428 78930
rect 57372 78866 57428 78878
rect 57820 78818 57876 78830
rect 57820 78766 57822 78818
rect 57874 78766 57876 78818
rect 57820 78596 57876 78766
rect 57820 78530 57876 78540
rect 56588 78094 56590 78146
rect 56642 78094 56644 78146
rect 55916 74834 55972 74844
rect 55244 74722 55300 74732
rect 54796 74174 54798 74226
rect 54850 74174 54852 74226
rect 54348 74162 54404 74172
rect 54796 74162 54852 74174
rect 52444 74062 52446 74114
rect 52498 74062 52500 74114
rect 52444 74050 52500 74062
rect 56364 74004 56420 76524
rect 56476 76356 56532 76366
rect 56476 76262 56532 76300
rect 56588 75796 56644 78094
rect 56700 78034 56756 78046
rect 56700 77982 56702 78034
rect 56754 77982 56756 78034
rect 56700 77924 56756 77982
rect 57820 78034 57876 78046
rect 57820 77982 57822 78034
rect 57874 77982 57876 78034
rect 56700 77858 56756 77868
rect 57372 77924 57428 77934
rect 57372 77830 57428 77868
rect 57484 77476 57540 77486
rect 57260 77474 57540 77476
rect 57260 77422 57486 77474
rect 57538 77422 57540 77474
rect 57260 77420 57540 77422
rect 57260 77362 57316 77420
rect 57484 77410 57540 77420
rect 57260 77310 57262 77362
rect 57314 77310 57316 77362
rect 57260 77298 57316 77310
rect 57708 77252 57764 77262
rect 57708 77158 57764 77196
rect 57372 77028 57428 77038
rect 57372 76356 57428 76972
rect 57596 76580 57652 76590
rect 57596 76486 57652 76524
rect 57708 76580 57764 76590
rect 57820 76580 57876 77982
rect 57708 76578 57876 76580
rect 57708 76526 57710 76578
rect 57762 76526 57876 76578
rect 57708 76524 57876 76526
rect 57708 76514 57764 76524
rect 57932 76356 57988 78932
rect 58268 78818 58324 78830
rect 58268 78766 58270 78818
rect 58322 78766 58324 78818
rect 58044 78146 58100 78158
rect 58044 78094 58046 78146
rect 58098 78094 58100 78146
rect 58044 78036 58100 78094
rect 58044 77970 58100 77980
rect 58156 78034 58212 78046
rect 58156 77982 58158 78034
rect 58210 77982 58212 78034
rect 58156 77924 58212 77982
rect 58156 77858 58212 77868
rect 58268 77476 58324 78766
rect 58380 78594 58436 78606
rect 58380 78542 58382 78594
rect 58434 78542 58436 78594
rect 58380 77700 58436 78542
rect 58380 77634 58436 77644
rect 58268 77474 58436 77476
rect 58268 77422 58270 77474
rect 58322 77422 58436 77474
rect 58268 77420 58436 77422
rect 58268 77410 58324 77420
rect 58156 77026 58212 77038
rect 58156 76974 58158 77026
rect 58210 76974 58212 77026
rect 58156 76580 58212 76974
rect 58156 76514 58212 76524
rect 58268 76692 58324 76702
rect 57932 76300 58212 76356
rect 56700 75796 56756 75806
rect 56588 75794 56756 75796
rect 56588 75742 56702 75794
rect 56754 75742 56756 75794
rect 56588 75740 56756 75742
rect 56700 75730 56756 75740
rect 57372 75682 57428 76300
rect 57596 76244 57652 76254
rect 57596 76242 58100 76244
rect 57596 76190 57598 76242
rect 57650 76190 58100 76242
rect 57596 76188 58100 76190
rect 57596 76178 57652 76188
rect 58044 75794 58100 76188
rect 58044 75742 58046 75794
rect 58098 75742 58100 75794
rect 58044 75730 58100 75742
rect 57372 75630 57374 75682
rect 57426 75630 57428 75682
rect 57372 75124 57428 75630
rect 57820 75124 57876 75134
rect 57372 75122 57876 75124
rect 57372 75070 57374 75122
rect 57426 75070 57822 75122
rect 57874 75070 57876 75122
rect 57372 75068 57876 75070
rect 57372 75058 57428 75068
rect 57820 75058 57876 75068
rect 56476 74788 56532 74798
rect 56476 74694 56532 74732
rect 57820 74004 57876 74014
rect 56364 73948 56532 74004
rect 51996 73892 52388 73948
rect 52332 73890 52388 73892
rect 52332 73838 52334 73890
rect 52386 73838 52388 73890
rect 50876 73218 51828 73220
rect 50876 73166 51326 73218
rect 51378 73166 51828 73218
rect 50876 73164 51828 73166
rect 51884 73220 51940 73230
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50428 71988 50484 71998
rect 50428 71894 50484 71932
rect 50764 71540 50820 71550
rect 50764 71446 50820 71484
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50316 69580 50484 69636
rect 50316 69300 50372 69310
rect 49980 69298 50372 69300
rect 49980 69246 50318 69298
rect 50370 69246 50372 69298
rect 49980 69244 50372 69246
rect 50316 69234 50372 69244
rect 50428 69076 50484 69580
rect 50316 69020 50484 69076
rect 50556 69020 50820 69030
rect 50204 68964 50260 68974
rect 50204 68850 50260 68908
rect 50204 68798 50206 68850
rect 50258 68798 50260 68850
rect 50204 68786 50260 68798
rect 49644 68628 49700 68638
rect 49644 67954 49700 68572
rect 49644 67902 49646 67954
rect 49698 67902 49700 67954
rect 49644 67890 49700 67902
rect 48972 67790 48974 67842
rect 49026 67790 49028 67842
rect 48972 67778 49028 67790
rect 50316 67284 50372 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 50540 68404 50596 68414
rect 50540 68310 50596 68348
rect 50988 68404 51044 68414
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 50204 67282 50372 67284
rect 50204 67230 50318 67282
rect 50370 67230 50372 67282
rect 50204 67228 50372 67230
rect 49756 67172 49812 67182
rect 49756 67078 49812 67116
rect 48860 67060 48916 67070
rect 48860 66966 48916 67004
rect 50092 67058 50148 67070
rect 50092 67006 50094 67058
rect 50146 67006 50148 67058
rect 48300 66948 48356 66958
rect 48300 66854 48356 66892
rect 49084 66948 49140 66958
rect 48860 64706 48916 64718
rect 48860 64654 48862 64706
rect 48914 64654 48916 64706
rect 48860 63812 48916 64654
rect 48860 63746 48916 63756
rect 48748 62468 48804 62478
rect 48748 62466 48916 62468
rect 48748 62414 48750 62466
rect 48802 62414 48916 62466
rect 48748 62412 48916 62414
rect 48748 62402 48804 62412
rect 48412 62354 48468 62366
rect 48412 62302 48414 62354
rect 48466 62302 48468 62354
rect 48412 61796 48468 62302
rect 47852 61740 48468 61796
rect 48860 62244 48916 62412
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 47628 60564 47684 60574
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 46956 59220 47012 59230
rect 46956 59126 47012 59164
rect 47628 59218 47684 60508
rect 47964 59444 48020 59454
rect 47852 59332 47908 59342
rect 47852 59238 47908 59276
rect 47628 59166 47630 59218
rect 47682 59166 47684 59218
rect 47628 59154 47684 59166
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 47964 58546 48020 59388
rect 47964 58494 47966 58546
rect 48018 58494 48020 58546
rect 47964 58482 48020 58494
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 2156 57092 2212 57102
rect 1820 37938 1876 37950
rect 1820 37886 1822 37938
rect 1874 37886 1876 37938
rect 1820 37492 1876 37886
rect 2156 37938 2212 57036
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 47964 54292 48020 54302
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 47964 53730 48020 54236
rect 47964 53678 47966 53730
rect 48018 53678 48020 53730
rect 47964 53666 48020 53678
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 48076 50036 48132 61740
rect 48860 61682 48916 62188
rect 48860 61630 48862 61682
rect 48914 61630 48916 61682
rect 48860 61618 48916 61630
rect 48412 60900 48468 60910
rect 48412 60806 48468 60844
rect 48748 60898 48804 60910
rect 48748 60846 48750 60898
rect 48802 60846 48804 60898
rect 48748 60340 48804 60846
rect 49084 60452 49140 66892
rect 49532 66276 49588 66286
rect 49532 66274 50036 66276
rect 49532 66222 49534 66274
rect 49586 66222 50036 66274
rect 49532 66220 50036 66222
rect 49532 66210 49588 66220
rect 49196 66162 49252 66174
rect 49196 66110 49198 66162
rect 49250 66110 49252 66162
rect 49196 65716 49252 66110
rect 49308 66052 49364 66062
rect 49868 66052 49924 66062
rect 49308 65958 49364 65996
rect 49644 66050 49924 66052
rect 49644 65998 49870 66050
rect 49922 65998 49924 66050
rect 49644 65996 49924 65998
rect 49644 65716 49700 65996
rect 49868 65986 49924 65996
rect 49196 65650 49252 65660
rect 49532 65660 49700 65716
rect 49980 65716 50036 66220
rect 50092 66162 50148 67006
rect 50204 66948 50260 67228
rect 50316 67218 50372 67228
rect 50428 67060 50484 67070
rect 50428 66966 50484 67004
rect 50988 66948 51044 68348
rect 51100 67620 51156 73164
rect 51324 73154 51380 73164
rect 51884 73126 51940 73164
rect 52332 73220 52388 73838
rect 56028 73442 56084 73454
rect 56028 73390 56030 73442
rect 56082 73390 56084 73442
rect 52332 73154 52388 73164
rect 53004 73220 53060 73230
rect 51548 71876 51604 71886
rect 51548 71874 51716 71876
rect 51548 71822 51550 71874
rect 51602 71822 51716 71874
rect 51548 71820 51716 71822
rect 51548 71810 51604 71820
rect 51436 71762 51492 71774
rect 51436 71710 51438 71762
rect 51490 71710 51492 71762
rect 51436 71652 51492 71710
rect 51436 71586 51492 71596
rect 51660 71090 51716 71820
rect 52108 71652 52164 71662
rect 52668 71652 52724 71662
rect 52108 71558 52164 71596
rect 52556 71650 52724 71652
rect 52556 71598 52670 71650
rect 52722 71598 52724 71650
rect 52556 71596 52724 71598
rect 51660 71038 51662 71090
rect 51714 71038 51716 71090
rect 51212 68852 51268 68862
rect 51212 68626 51268 68796
rect 51324 68740 51380 68750
rect 51660 68740 51716 71038
rect 52556 71540 52612 71596
rect 52668 71586 52724 71596
rect 52780 71652 52836 71662
rect 52108 70754 52164 70766
rect 52108 70702 52110 70754
rect 52162 70702 52164 70754
rect 52108 70532 52164 70702
rect 52108 70466 52164 70476
rect 52444 69524 52500 69534
rect 52556 69524 52612 71484
rect 52444 69522 52612 69524
rect 52444 69470 52446 69522
rect 52498 69470 52612 69522
rect 52444 69468 52612 69470
rect 52668 70754 52724 70766
rect 52668 70702 52670 70754
rect 52722 70702 52724 70754
rect 52668 70532 52724 70702
rect 51324 68738 51716 68740
rect 51324 68686 51326 68738
rect 51378 68686 51716 68738
rect 51324 68684 51716 68686
rect 52108 68738 52164 68750
rect 52108 68686 52110 68738
rect 52162 68686 52164 68738
rect 51324 68674 51380 68684
rect 51212 68574 51214 68626
rect 51266 68574 51268 68626
rect 51212 68562 51268 68574
rect 51884 68628 51940 68638
rect 51884 68534 51940 68572
rect 52108 68066 52164 68686
rect 52220 68628 52276 68638
rect 52220 68626 52388 68628
rect 52220 68574 52222 68626
rect 52274 68574 52388 68626
rect 52220 68572 52388 68574
rect 52220 68562 52276 68572
rect 52108 68014 52110 68066
rect 52162 68014 52164 68066
rect 52108 68002 52164 68014
rect 51772 67956 51828 67966
rect 51772 67954 52052 67956
rect 51772 67902 51774 67954
rect 51826 67902 52052 67954
rect 51772 67900 52052 67902
rect 51772 67890 51828 67900
rect 51100 67554 51156 67564
rect 51996 67282 52052 67900
rect 51996 67230 51998 67282
rect 52050 67230 52052 67282
rect 51996 67218 52052 67230
rect 52108 67620 52164 67630
rect 52220 67620 52276 67630
rect 52164 67618 52276 67620
rect 52164 67566 52222 67618
rect 52274 67566 52276 67618
rect 52164 67564 52276 67566
rect 51100 67172 51156 67182
rect 51100 67078 51156 67116
rect 51212 67172 51268 67182
rect 51884 67172 51940 67182
rect 51212 67170 51380 67172
rect 51212 67118 51214 67170
rect 51266 67118 51380 67170
rect 51212 67116 51380 67118
rect 51212 67106 51268 67116
rect 50988 66892 51156 66948
rect 50204 66882 50260 66892
rect 50092 66110 50094 66162
rect 50146 66110 50148 66162
rect 50092 66098 50148 66110
rect 50204 66164 50260 66174
rect 50204 66070 50260 66108
rect 50988 66162 51044 66174
rect 50988 66110 50990 66162
rect 51042 66110 51044 66162
rect 50652 66052 50708 66062
rect 50428 66050 50708 66052
rect 50428 65998 50654 66050
rect 50706 65998 50708 66050
rect 50428 65996 50708 65998
rect 49980 65660 50372 65716
rect 49532 64818 49588 65660
rect 50316 65602 50372 65660
rect 50316 65550 50318 65602
rect 50370 65550 50372 65602
rect 50316 65538 50372 65550
rect 49532 64766 49534 64818
rect 49586 64766 49588 64818
rect 49532 64754 49588 64766
rect 49644 65490 49700 65502
rect 49644 65438 49646 65490
rect 49698 65438 49700 65490
rect 49532 63924 49588 63934
rect 49644 63924 49700 65438
rect 50428 64596 50484 65996
rect 50652 65986 50708 65996
rect 50876 66050 50932 66062
rect 50876 65998 50878 66050
rect 50930 65998 50932 66050
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 50876 65716 50932 65998
rect 50876 65650 50932 65660
rect 49532 63922 49700 63924
rect 49532 63870 49534 63922
rect 49586 63870 49700 63922
rect 49532 63868 49700 63870
rect 50092 64540 50484 64596
rect 50540 65604 50596 65614
rect 49532 63812 49588 63868
rect 49420 63140 49476 63150
rect 49532 63140 49588 63756
rect 50092 63250 50148 64540
rect 50540 64484 50596 65548
rect 50988 64708 51044 66110
rect 50988 64642 51044 64652
rect 50316 64428 50596 64484
rect 50316 64034 50372 64428
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 50316 63982 50318 64034
rect 50370 63982 50372 64034
rect 50316 63970 50372 63982
rect 50092 63198 50094 63250
rect 50146 63198 50148 63250
rect 50092 63186 50148 63198
rect 50316 63476 50372 63486
rect 49420 63138 49588 63140
rect 49420 63086 49422 63138
rect 49474 63086 49588 63138
rect 49420 63084 49588 63086
rect 49420 62916 49476 63084
rect 49420 62850 49476 62860
rect 50316 62244 50372 63420
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 49756 61572 49812 61582
rect 49756 61570 49924 61572
rect 49756 61518 49758 61570
rect 49810 61518 49924 61570
rect 49756 61516 49924 61518
rect 49756 61506 49812 61516
rect 49420 61346 49476 61358
rect 49420 61294 49422 61346
rect 49474 61294 49476 61346
rect 49420 60900 49476 61294
rect 49420 60834 49476 60844
rect 49868 60788 49924 61516
rect 50316 61458 50372 62188
rect 51100 62188 51156 66892
rect 51324 64820 51380 67116
rect 51884 67078 51940 67116
rect 51436 67060 51492 67070
rect 51436 67058 51716 67060
rect 51436 67006 51438 67058
rect 51490 67006 51716 67058
rect 51436 67004 51716 67006
rect 51436 66994 51492 67004
rect 51660 66164 51716 67004
rect 51436 66050 51492 66062
rect 51436 65998 51438 66050
rect 51490 65998 51492 66050
rect 51660 66032 51716 66108
rect 51772 66164 51828 66174
rect 51772 66162 52052 66164
rect 51772 66110 51774 66162
rect 51826 66110 52052 66162
rect 51772 66108 52052 66110
rect 51772 66098 51828 66108
rect 51436 65604 51492 65998
rect 51436 65538 51492 65548
rect 51772 65828 51828 65838
rect 51660 64820 51716 64830
rect 51324 64818 51716 64820
rect 51324 64766 51662 64818
rect 51714 64766 51716 64818
rect 51324 64764 51716 64766
rect 51660 64754 51716 64764
rect 51772 64596 51828 65772
rect 51996 64708 52052 66108
rect 52108 65828 52164 67564
rect 52220 67554 52276 67564
rect 52220 67060 52276 67070
rect 52332 67060 52388 68572
rect 52444 68402 52500 69468
rect 52668 69412 52724 70476
rect 52668 69188 52724 69356
rect 52668 68850 52724 69132
rect 52668 68798 52670 68850
rect 52722 68798 52724 68850
rect 52668 68786 52724 68798
rect 52780 68852 52836 71596
rect 52892 70196 52948 70206
rect 52892 70102 52948 70140
rect 52780 68786 52836 68796
rect 53004 68628 53060 73164
rect 53900 72548 53956 72558
rect 53788 71762 53844 71774
rect 53788 71710 53790 71762
rect 53842 71710 53844 71762
rect 53340 71650 53396 71662
rect 53340 71598 53342 71650
rect 53394 71598 53396 71650
rect 53340 70756 53396 71598
rect 53340 70690 53396 70700
rect 53564 70866 53620 70878
rect 53564 70814 53566 70866
rect 53618 70814 53620 70866
rect 53564 70756 53620 70814
rect 53564 70690 53620 70700
rect 53676 70532 53732 70542
rect 53788 70532 53844 71710
rect 53900 70866 53956 72492
rect 55468 72436 55524 72446
rect 55468 72342 55524 72380
rect 54684 72324 54740 72334
rect 55132 72324 55188 72334
rect 54684 72230 54740 72268
rect 54796 72322 55188 72324
rect 54796 72270 55134 72322
rect 55186 72270 55188 72322
rect 54796 72268 55188 72270
rect 54796 71988 54852 72268
rect 55132 72258 55188 72268
rect 55244 72324 55300 72334
rect 54572 71932 54852 71988
rect 54572 71874 54628 71932
rect 54572 71822 54574 71874
rect 54626 71822 54628 71874
rect 54572 71810 54628 71822
rect 53900 70814 53902 70866
rect 53954 70814 53956 70866
rect 53900 70802 53956 70814
rect 55132 70978 55188 70990
rect 55132 70926 55134 70978
rect 55186 70926 55188 70978
rect 53732 70476 53844 70532
rect 55132 70532 55188 70926
rect 53676 69410 53732 70476
rect 55132 70466 55188 70476
rect 53676 69358 53678 69410
rect 53730 69358 53732 69410
rect 53676 69188 53732 69358
rect 54572 69972 54628 69982
rect 52444 68350 52446 68402
rect 52498 68350 52500 68402
rect 52444 68338 52500 68350
rect 52780 68572 53060 68628
rect 53564 69132 53676 69188
rect 52556 68066 52612 68078
rect 52556 68014 52558 68066
rect 52610 68014 52612 68066
rect 52556 67282 52612 68014
rect 52668 67620 52724 67630
rect 52780 67620 52836 68572
rect 53116 68514 53172 68526
rect 53116 68462 53118 68514
rect 53170 68462 53172 68514
rect 53004 68402 53060 68414
rect 53004 68350 53006 68402
rect 53058 68350 53060 68402
rect 52668 67618 52836 67620
rect 52668 67566 52670 67618
rect 52722 67566 52836 67618
rect 52668 67564 52836 67566
rect 52668 67554 52724 67564
rect 52556 67230 52558 67282
rect 52610 67230 52612 67282
rect 52556 67218 52612 67230
rect 52780 67282 52836 67564
rect 52780 67230 52782 67282
rect 52834 67230 52836 67282
rect 52220 67058 52388 67060
rect 52220 67006 52222 67058
rect 52274 67006 52388 67058
rect 52220 67004 52388 67006
rect 52220 66994 52276 67004
rect 52220 66052 52276 66062
rect 52220 65958 52276 65996
rect 52332 65940 52388 67004
rect 52556 66276 52612 66286
rect 52556 66182 52612 66220
rect 52332 65874 52388 65884
rect 52444 66050 52500 66062
rect 52444 65998 52446 66050
rect 52498 65998 52500 66050
rect 52108 65762 52164 65772
rect 52444 65828 52500 65998
rect 52444 65762 52500 65772
rect 52444 65604 52500 65614
rect 52444 65378 52500 65548
rect 52444 65326 52446 65378
rect 52498 65326 52500 65378
rect 52444 65314 52500 65326
rect 52108 64708 52164 64718
rect 51996 64706 52164 64708
rect 51996 64654 52110 64706
rect 52162 64654 52164 64706
rect 51996 64652 52164 64654
rect 52108 64642 52164 64652
rect 51660 64540 51828 64596
rect 52444 64596 52500 64606
rect 51100 62132 51380 62188
rect 50316 61406 50318 61458
rect 50370 61406 50372 61458
rect 50316 61394 50372 61406
rect 50428 61570 50484 61582
rect 50428 61518 50430 61570
rect 50482 61518 50484 61570
rect 50092 60788 50148 60798
rect 49868 60786 50148 60788
rect 49868 60734 50094 60786
rect 50146 60734 50148 60786
rect 49868 60732 50148 60734
rect 49756 60564 49812 60574
rect 49756 60470 49812 60508
rect 49084 60396 49252 60452
rect 48748 60284 49140 60340
rect 49084 60114 49140 60284
rect 49084 60062 49086 60114
rect 49138 60062 49140 60114
rect 49084 60050 49140 60062
rect 48412 60004 48468 60014
rect 48412 59910 48468 59948
rect 48748 59444 48804 59454
rect 48748 59350 48804 59388
rect 49196 59444 49252 60396
rect 50092 60116 50148 60732
rect 50428 60788 50484 61518
rect 51100 61346 51156 61358
rect 51100 61294 51102 61346
rect 51154 61294 51156 61346
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50876 60898 50932 60910
rect 50876 60846 50878 60898
rect 50930 60846 50932 60898
rect 50428 60722 50484 60732
rect 50764 60788 50820 60798
rect 50764 60694 50820 60732
rect 50876 60676 50932 60846
rect 51100 60788 51156 61294
rect 51100 60722 51156 60732
rect 50876 60610 50932 60620
rect 50092 60050 50148 60060
rect 51212 60116 51268 60126
rect 51212 60022 51268 60060
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 49196 59378 49252 59388
rect 50428 59444 50484 59454
rect 50316 59332 50372 59342
rect 50316 59238 50372 59276
rect 48524 59220 48580 59230
rect 48524 59126 48580 59164
rect 49532 59218 49588 59230
rect 49532 59166 49534 59218
rect 49586 59166 49588 59218
rect 48524 58436 48580 58446
rect 48524 58342 48580 58380
rect 49420 58436 49476 58446
rect 49420 58342 49476 58380
rect 48748 58212 48804 58222
rect 48748 58210 49140 58212
rect 48748 58158 48750 58210
rect 48802 58158 49140 58210
rect 48748 58156 49140 58158
rect 48748 58146 48804 58156
rect 49084 56978 49140 58156
rect 49084 56926 49086 56978
rect 49138 56926 49140 56978
rect 49084 56914 49140 56926
rect 48412 56866 48468 56878
rect 48412 56814 48414 56866
rect 48466 56814 48468 56866
rect 48300 56420 48356 56430
rect 48300 54628 48356 56364
rect 48412 56308 48468 56814
rect 48412 55300 48468 56252
rect 49532 56308 49588 59166
rect 49756 58434 49812 58446
rect 49756 58382 49758 58434
rect 49810 58382 49812 58434
rect 49644 57426 49700 57438
rect 49644 57374 49646 57426
rect 49698 57374 49700 57426
rect 49644 56420 49700 57374
rect 49756 56980 49812 58382
rect 50428 58322 50484 59388
rect 51100 58658 51156 58670
rect 51100 58606 51102 58658
rect 51154 58606 51156 58658
rect 50540 58548 50596 58558
rect 51100 58548 51156 58606
rect 50540 58434 50596 58492
rect 50540 58382 50542 58434
rect 50594 58382 50596 58434
rect 50540 58370 50596 58382
rect 50876 58546 51156 58548
rect 50876 58494 51102 58546
rect 51154 58494 51156 58546
rect 50876 58492 51156 58494
rect 50428 58270 50430 58322
rect 50482 58270 50484 58322
rect 50428 58258 50484 58270
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50876 57876 50932 58492
rect 50652 57820 50932 57876
rect 50652 57762 50708 57820
rect 50652 57710 50654 57762
rect 50706 57710 50708 57762
rect 50652 57698 50708 57710
rect 50764 57650 50820 57662
rect 50764 57598 50766 57650
rect 50818 57598 50820 57650
rect 50764 57540 50820 57598
rect 50764 57474 50820 57484
rect 49756 56914 49812 56924
rect 49980 57426 50036 57438
rect 49980 57374 49982 57426
rect 50034 57374 50036 57426
rect 49644 56354 49700 56364
rect 49532 56242 49588 56252
rect 49980 55468 50036 57374
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 50652 56308 50708 56318
rect 50652 56214 50708 56252
rect 49980 55412 50260 55468
rect 48412 55298 48580 55300
rect 48412 55246 48414 55298
rect 48466 55246 48580 55298
rect 48412 55244 48580 55246
rect 48412 55234 48468 55244
rect 48412 54628 48468 54638
rect 48300 54626 48468 54628
rect 48300 54574 48414 54626
rect 48466 54574 48468 54626
rect 48300 54572 48468 54574
rect 48412 54562 48468 54572
rect 48524 54516 48580 55244
rect 49084 55186 49140 55198
rect 49084 55134 49086 55186
rect 49138 55134 49140 55186
rect 48748 54738 48804 54750
rect 48748 54686 48750 54738
rect 48802 54686 48804 54738
rect 48748 54628 48804 54686
rect 49084 54628 49140 55134
rect 48748 54572 49140 54628
rect 48524 54460 48916 54516
rect 48860 53730 48916 54460
rect 50204 54514 50260 55356
rect 51100 55188 51156 58492
rect 51324 57876 51380 62132
rect 51436 60676 51492 60686
rect 51436 60582 51492 60620
rect 51660 58658 51716 64540
rect 52444 64502 52500 64540
rect 52332 64482 52388 64494
rect 52332 64430 52334 64482
rect 52386 64430 52388 64482
rect 52332 63924 52388 64430
rect 52444 63924 52500 63934
rect 52332 63868 52444 63924
rect 52444 63810 52500 63868
rect 52444 63758 52446 63810
rect 52498 63758 52500 63810
rect 52444 63746 52500 63758
rect 52780 63476 52836 67230
rect 52892 67620 52948 67630
rect 52892 67170 52948 67564
rect 52892 67118 52894 67170
rect 52946 67118 52948 67170
rect 52892 67060 52948 67118
rect 52892 66276 52948 67004
rect 52892 66210 52948 66220
rect 52892 63924 52948 63934
rect 53004 63924 53060 68350
rect 53116 68404 53172 68462
rect 53116 68338 53172 68348
rect 53340 67620 53396 67630
rect 53340 67526 53396 67564
rect 53228 67172 53284 67182
rect 53116 65604 53172 65614
rect 53116 65510 53172 65548
rect 53228 65602 53284 67116
rect 53452 66946 53508 66958
rect 53452 66894 53454 66946
rect 53506 66894 53508 66946
rect 53228 65550 53230 65602
rect 53282 65550 53284 65602
rect 53228 65538 53284 65550
rect 53340 65716 53396 65726
rect 53116 65268 53172 65278
rect 53340 65268 53396 65660
rect 53116 65266 53396 65268
rect 53116 65214 53118 65266
rect 53170 65214 53396 65266
rect 53116 65212 53396 65214
rect 53116 65202 53172 65212
rect 53452 64932 53508 66894
rect 53564 66274 53620 69132
rect 53676 69122 53732 69132
rect 54348 69298 54404 69310
rect 54348 69246 54350 69298
rect 54402 69246 54404 69298
rect 53676 68852 53732 68862
rect 53676 68758 53732 68796
rect 54236 68852 54292 68862
rect 54348 68852 54404 69246
rect 54236 68850 54404 68852
rect 54236 68798 54238 68850
rect 54290 68798 54404 68850
rect 54236 68796 54404 68798
rect 54236 68786 54292 68796
rect 54572 68738 54628 69916
rect 55132 68852 55188 68862
rect 55244 68852 55300 72268
rect 56028 72100 56084 73390
rect 56364 73330 56420 73342
rect 56364 73278 56366 73330
rect 56418 73278 56420 73330
rect 56364 72772 56420 73278
rect 56364 72706 56420 72716
rect 56476 73220 56532 73948
rect 56476 72546 56532 73164
rect 56476 72494 56478 72546
rect 56530 72494 56532 72546
rect 56140 72436 56196 72446
rect 56140 72342 56196 72380
rect 56476 72324 56532 72494
rect 57148 73892 57204 73902
rect 57148 72546 57204 73836
rect 57484 73220 57540 73230
rect 57148 72494 57150 72546
rect 57202 72494 57204 72546
rect 57148 72482 57204 72494
rect 57372 73218 57540 73220
rect 57372 73166 57486 73218
rect 57538 73166 57540 73218
rect 57372 73164 57540 73166
rect 56476 72258 56532 72268
rect 57260 72434 57316 72446
rect 57260 72382 57262 72434
rect 57314 72382 57316 72434
rect 55804 72044 56084 72100
rect 55804 71090 55860 72044
rect 56700 71652 56756 71662
rect 56700 71558 56756 71596
rect 57260 71652 57316 72382
rect 57260 71586 57316 71596
rect 55804 71038 55806 71090
rect 55858 71038 55860 71090
rect 55804 71026 55860 71038
rect 57372 70644 57428 73164
rect 57484 73154 57540 73164
rect 57820 73218 57876 73948
rect 58156 74004 58212 76300
rect 58268 76244 58324 76636
rect 58380 76690 58436 77420
rect 58380 76638 58382 76690
rect 58434 76638 58436 76690
rect 58380 76626 58436 76638
rect 58492 76692 58548 79662
rect 58828 78932 58884 78942
rect 58828 78706 58884 78876
rect 58940 78820 58996 81902
rect 59500 81842 59556 85148
rect 60284 85202 60340 87836
rect 60508 87332 60564 87948
rect 60620 87938 60676 87948
rect 61516 88002 61572 88014
rect 61516 87950 61518 88002
rect 61570 87950 61572 88002
rect 60284 85150 60286 85202
rect 60338 85150 60340 85202
rect 60396 85762 60452 85774
rect 60396 85710 60398 85762
rect 60450 85710 60452 85762
rect 60396 85316 60452 85710
rect 60508 85764 60564 87276
rect 60620 87332 60676 87342
rect 60620 87330 61460 87332
rect 60620 87278 60622 87330
rect 60674 87278 61460 87330
rect 60620 87276 61460 87278
rect 60620 87266 60676 87276
rect 60844 86996 60900 87006
rect 60508 85698 60564 85708
rect 60620 86772 60676 86782
rect 60452 85260 60564 85316
rect 60396 85184 60452 85260
rect 60284 85138 60340 85150
rect 60396 82628 60452 82638
rect 60396 82534 60452 82572
rect 59500 81790 59502 81842
rect 59554 81790 59556 81842
rect 59500 81778 59556 81790
rect 59724 81954 59780 81966
rect 59724 81902 59726 81954
rect 59778 81902 59780 81954
rect 59724 81732 59780 81902
rect 59724 81666 59780 81676
rect 60284 81732 60340 81742
rect 60284 81638 60340 81676
rect 59500 79828 59556 79838
rect 59052 79602 59108 79614
rect 59052 79550 59054 79602
rect 59106 79550 59108 79602
rect 59052 79044 59108 79550
rect 59500 79602 59556 79772
rect 59500 79550 59502 79602
rect 59554 79550 59556 79602
rect 59500 79538 59556 79550
rect 60508 79602 60564 85260
rect 60620 84420 60676 86716
rect 60844 85540 60900 86940
rect 61404 86546 61460 87276
rect 61516 86660 61572 87950
rect 61852 87332 61908 88174
rect 62524 88226 62580 88238
rect 62524 88174 62526 88226
rect 62578 88174 62580 88226
rect 62524 87892 62580 88174
rect 62636 88116 62692 88126
rect 62636 88114 62804 88116
rect 62636 88062 62638 88114
rect 62690 88062 62804 88114
rect 62636 88060 62804 88062
rect 62636 88050 62692 88060
rect 62524 87826 62580 87836
rect 61852 87266 61908 87276
rect 62748 87556 62804 88060
rect 62748 87330 62804 87500
rect 62748 87278 62750 87330
rect 62802 87278 62804 87330
rect 62748 87266 62804 87278
rect 62412 87220 62468 87230
rect 62188 86772 62244 86782
rect 62188 86678 62244 86716
rect 61628 86660 61684 86670
rect 61516 86658 61684 86660
rect 61516 86606 61630 86658
rect 61682 86606 61684 86658
rect 61516 86604 61684 86606
rect 61628 86594 61684 86604
rect 61404 86494 61406 86546
rect 61458 86494 61460 86546
rect 61404 86482 61460 86494
rect 61516 86212 61572 86222
rect 60956 85764 61012 85774
rect 60956 85670 61012 85708
rect 60844 85484 61012 85540
rect 60620 84418 60900 84420
rect 60620 84366 60622 84418
rect 60674 84366 60900 84418
rect 60620 84364 60900 84366
rect 60620 84354 60676 84364
rect 60844 82962 60900 84364
rect 60844 82910 60846 82962
rect 60898 82910 60900 82962
rect 60844 82068 60900 82910
rect 60620 82012 60844 82068
rect 60620 81170 60676 82012
rect 60844 82002 60900 82012
rect 60620 81118 60622 81170
rect 60674 81118 60676 81170
rect 60620 81106 60676 81118
rect 60508 79550 60510 79602
rect 60562 79550 60564 79602
rect 60508 79538 60564 79550
rect 59052 78978 59108 78988
rect 59500 79380 59556 79390
rect 59388 78820 59444 78830
rect 58940 78818 59444 78820
rect 58940 78766 59390 78818
rect 59442 78766 59444 78818
rect 58940 78764 59444 78766
rect 59388 78754 59444 78764
rect 58828 78654 58830 78706
rect 58882 78654 58884 78706
rect 58828 78372 58884 78654
rect 58828 78306 58884 78316
rect 59276 78148 59332 78158
rect 59500 78148 59556 79324
rect 60956 78988 61012 85484
rect 61516 85090 61572 86156
rect 61516 85038 61518 85090
rect 61570 85038 61572 85090
rect 61516 85026 61572 85038
rect 61740 85876 61796 85886
rect 61740 84978 61796 85820
rect 61740 84926 61742 84978
rect 61794 84926 61796 84978
rect 61740 84914 61796 84926
rect 62412 85764 62468 87164
rect 63084 87220 63140 88846
rect 63084 87154 63140 87164
rect 63308 88898 63588 88900
rect 63308 88846 63534 88898
rect 63586 88846 63588 88898
rect 63308 88844 63588 88846
rect 63308 86772 63364 88844
rect 63532 88834 63588 88844
rect 65916 88620 66180 88630
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 65916 88554 66180 88564
rect 63532 88114 63588 88126
rect 63532 88062 63534 88114
rect 63586 88062 63588 88114
rect 63308 86706 63364 86716
rect 63420 87218 63476 87230
rect 63420 87166 63422 87218
rect 63474 87166 63476 87218
rect 61628 82852 61684 82862
rect 61292 82850 61684 82852
rect 61292 82798 61630 82850
rect 61682 82798 61684 82850
rect 61292 82796 61684 82798
rect 61292 81282 61348 82796
rect 61628 82786 61684 82796
rect 61964 82740 62020 82750
rect 61964 82738 62132 82740
rect 61964 82686 61966 82738
rect 62018 82686 62132 82738
rect 61964 82684 62132 82686
rect 61964 82674 62020 82684
rect 62076 82180 62132 82684
rect 62300 82180 62356 82190
rect 62076 82178 62356 82180
rect 62076 82126 62302 82178
rect 62354 82126 62356 82178
rect 62076 82124 62356 82126
rect 62300 82114 62356 82124
rect 61292 81230 61294 81282
rect 61346 81230 61348 81282
rect 61292 81218 61348 81230
rect 62188 81956 62244 81966
rect 61516 80612 61572 80622
rect 61404 80500 61460 80510
rect 61404 80406 61460 80444
rect 61180 79492 61236 79502
rect 61180 79398 61236 79436
rect 60508 78932 61012 78988
rect 60396 78820 60452 78830
rect 60396 78726 60452 78764
rect 59276 78146 59556 78148
rect 59276 78094 59278 78146
rect 59330 78094 59556 78146
rect 59276 78092 59556 78094
rect 59724 78596 59780 78606
rect 59276 78082 59332 78092
rect 59724 78034 59780 78540
rect 60284 78146 60340 78158
rect 60284 78094 60286 78146
rect 60338 78094 60340 78146
rect 59724 77982 59726 78034
rect 59778 77982 59780 78034
rect 59724 77970 59780 77982
rect 60060 78036 60116 78046
rect 60116 77980 60228 78036
rect 60060 77942 60116 77980
rect 58604 77924 58660 77934
rect 58660 77868 58772 77924
rect 58604 77792 58660 77868
rect 58604 77028 58660 77038
rect 58716 77028 58772 77868
rect 58940 77028 58996 77038
rect 58716 76972 58940 77028
rect 58604 76934 58660 76972
rect 58492 76636 58660 76692
rect 58492 76468 58548 76478
rect 58492 76374 58548 76412
rect 58380 76244 58436 76254
rect 58268 76242 58436 76244
rect 58268 76190 58382 76242
rect 58434 76190 58436 76242
rect 58268 76188 58436 76190
rect 58380 76178 58436 76188
rect 58604 73948 58660 76636
rect 58940 76690 58996 76972
rect 58940 76638 58942 76690
rect 58994 76638 58996 76690
rect 58940 76468 58996 76638
rect 58940 76402 58996 76412
rect 60172 75794 60228 77980
rect 60172 75742 60174 75794
rect 60226 75742 60228 75794
rect 60172 75730 60228 75742
rect 58156 73938 58212 73948
rect 58268 73892 58324 73902
rect 58268 73554 58324 73836
rect 58268 73502 58270 73554
rect 58322 73502 58324 73554
rect 58268 73490 58324 73502
rect 58492 73892 58660 73948
rect 59724 74004 59780 74014
rect 60284 73948 60340 78094
rect 60396 74116 60452 74126
rect 60396 74022 60452 74060
rect 59724 73910 59780 73948
rect 59500 73892 59556 73902
rect 57820 73166 57822 73218
rect 57874 73166 57876 73218
rect 57820 72548 57876 73166
rect 58044 72772 58100 72782
rect 58044 72678 58100 72716
rect 57820 72482 57876 72492
rect 58380 72548 58436 72558
rect 58380 72454 58436 72492
rect 58492 71876 58548 73892
rect 59500 73554 59556 73836
rect 59500 73502 59502 73554
rect 59554 73502 59556 73554
rect 59500 72660 59556 73502
rect 59836 73892 60340 73948
rect 59724 72660 59780 72670
rect 59164 72658 59780 72660
rect 59164 72606 59726 72658
rect 59778 72606 59780 72658
rect 59164 72604 59780 72606
rect 59164 72546 59220 72604
rect 59724 72594 59780 72604
rect 59164 72494 59166 72546
rect 59218 72494 59220 72546
rect 58268 71820 58548 71876
rect 59052 72434 59108 72446
rect 59052 72382 59054 72434
rect 59106 72382 59108 72434
rect 57932 71092 57988 71102
rect 57932 70998 57988 71036
rect 56476 70532 56532 70542
rect 56252 70420 56308 70430
rect 55132 68850 55300 68852
rect 55132 68798 55134 68850
rect 55186 68798 55300 68850
rect 55132 68796 55300 68798
rect 55580 70196 55636 70206
rect 55132 68786 55188 68796
rect 54572 68686 54574 68738
rect 54626 68686 54628 68738
rect 54572 68674 54628 68686
rect 54684 68740 54740 68750
rect 53788 67620 53844 67630
rect 53788 67526 53844 67564
rect 54236 67508 54292 67518
rect 53788 67172 53844 67182
rect 54236 67172 54292 67452
rect 53844 67170 54292 67172
rect 53844 67118 54238 67170
rect 54290 67118 54292 67170
rect 53844 67116 54292 67118
rect 53788 67040 53844 67116
rect 54236 67106 54292 67116
rect 54684 66836 54740 68684
rect 55356 68626 55412 68638
rect 55356 68574 55358 68626
rect 55410 68574 55412 68626
rect 54796 67620 54852 67630
rect 55356 67620 55412 68574
rect 54796 67618 55412 67620
rect 54796 67566 54798 67618
rect 54850 67566 55412 67618
rect 54796 67564 55412 67566
rect 54796 67554 54852 67564
rect 54684 66770 54740 66780
rect 53564 66222 53566 66274
rect 53618 66222 53620 66274
rect 53564 66210 53620 66222
rect 54348 66164 54404 66174
rect 53788 66162 54404 66164
rect 53788 66110 54350 66162
rect 54402 66110 54404 66162
rect 53788 66108 54404 66110
rect 53788 65714 53844 66108
rect 54348 66098 54404 66108
rect 53788 65662 53790 65714
rect 53842 65662 53844 65714
rect 53788 65650 53844 65662
rect 54012 65940 54068 65950
rect 54012 65714 54068 65884
rect 54012 65662 54014 65714
rect 54066 65662 54068 65714
rect 54012 65650 54068 65662
rect 54124 65604 54180 65614
rect 54124 65510 54180 65548
rect 54572 65492 54628 65502
rect 54572 65398 54628 65436
rect 53340 64708 53396 64718
rect 53340 64614 53396 64652
rect 53452 64036 53508 64876
rect 53676 65268 53732 65278
rect 53676 64706 53732 65212
rect 54124 64932 54180 64942
rect 54124 64820 54180 64876
rect 54572 64820 54628 64830
rect 54124 64818 54628 64820
rect 54124 64766 54126 64818
rect 54178 64766 54574 64818
rect 54626 64766 54628 64818
rect 54124 64764 54628 64766
rect 54124 64754 54180 64764
rect 54572 64754 54628 64764
rect 53676 64654 53678 64706
rect 53730 64654 53732 64706
rect 53676 64596 53732 64654
rect 53676 64530 53732 64540
rect 54684 64596 54740 64606
rect 52892 63922 53060 63924
rect 52892 63870 52894 63922
rect 52946 63870 53060 63922
rect 52892 63868 53060 63870
rect 53340 63980 53508 64036
rect 53564 64482 53620 64494
rect 53564 64430 53566 64482
rect 53618 64430 53620 64482
rect 52892 63476 52948 63868
rect 53004 63476 53060 63486
rect 52892 63420 53004 63476
rect 52780 63410 52836 63420
rect 53004 63410 53060 63420
rect 52220 63250 52276 63262
rect 52220 63198 52222 63250
rect 52274 63198 52276 63250
rect 52220 63140 52276 63198
rect 52220 63074 52276 63084
rect 52668 63252 52724 63262
rect 51772 62916 51828 62926
rect 51772 62468 51828 62860
rect 51772 60004 51828 62412
rect 52668 62468 52724 63196
rect 53340 63252 53396 63980
rect 53340 63186 53396 63196
rect 53452 63812 53508 63822
rect 52668 62336 52724 62412
rect 53452 62188 53508 63756
rect 53564 63140 53620 64430
rect 54460 64034 54516 64046
rect 54460 63982 54462 64034
rect 54514 63982 54516 64034
rect 53900 63922 53956 63934
rect 53900 63870 53902 63922
rect 53954 63870 53956 63922
rect 53900 63140 53956 63870
rect 54236 63924 54292 63934
rect 54236 63830 54292 63868
rect 54460 63364 54516 63982
rect 54460 63298 54516 63308
rect 54124 63140 54180 63150
rect 53900 63138 54180 63140
rect 53900 63086 54126 63138
rect 54178 63086 54180 63138
rect 53900 63084 54180 63086
rect 53564 63074 53620 63084
rect 53228 62132 53508 62188
rect 53676 63026 53732 63038
rect 53676 62974 53678 63026
rect 53730 62974 53732 63026
rect 52332 61348 52388 61358
rect 51884 60788 51940 60798
rect 51884 60676 51940 60732
rect 51884 60674 52052 60676
rect 51884 60622 51886 60674
rect 51938 60622 52052 60674
rect 51884 60620 52052 60622
rect 51884 60610 51940 60620
rect 51772 59910 51828 59948
rect 51660 58606 51662 58658
rect 51714 58606 51716 58658
rect 51660 58594 51716 58606
rect 51996 58548 52052 60620
rect 51996 58454 52052 58492
rect 51660 58212 51716 58222
rect 51660 58210 51828 58212
rect 51660 58158 51662 58210
rect 51714 58158 51828 58210
rect 51660 58156 51828 58158
rect 51660 58146 51716 58156
rect 51436 57876 51492 57886
rect 51324 57874 51492 57876
rect 51324 57822 51438 57874
rect 51490 57822 51492 57874
rect 51324 57820 51492 57822
rect 51436 57810 51492 57820
rect 51772 57652 51828 58156
rect 51772 57650 52164 57652
rect 51772 57598 51774 57650
rect 51826 57598 52164 57650
rect 51772 57596 52164 57598
rect 51772 57586 51828 57596
rect 51212 56980 51268 56990
rect 51212 56886 51268 56924
rect 51996 56980 52052 56990
rect 51660 56644 51716 56654
rect 51436 56642 51716 56644
rect 51436 56590 51662 56642
rect 51714 56590 51716 56642
rect 51436 56588 51716 56590
rect 51436 56308 51492 56588
rect 51660 56578 51716 56588
rect 51436 56194 51492 56252
rect 51436 56142 51438 56194
rect 51490 56142 51492 56194
rect 51436 56130 51492 56142
rect 51212 55412 51268 55422
rect 51212 55318 51268 55356
rect 51772 55188 51828 55198
rect 51100 55186 51828 55188
rect 51100 55134 51774 55186
rect 51826 55134 51828 55186
rect 51100 55132 51828 55134
rect 51772 55122 51828 55132
rect 51996 54964 52052 56924
rect 52108 55188 52164 57596
rect 52220 57540 52276 57550
rect 52220 57446 52276 57484
rect 52108 55094 52164 55132
rect 52220 56308 52276 56318
rect 50556 54908 50820 54918
rect 51996 54908 52164 54964
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50204 54462 50206 54514
rect 50258 54462 50260 54514
rect 50204 54450 50260 54462
rect 50876 54626 50932 54638
rect 50876 54574 50878 54626
rect 50930 54574 50932 54626
rect 49868 54292 49924 54302
rect 48860 53678 48862 53730
rect 48914 53678 48916 53730
rect 48188 53620 48244 53630
rect 48188 53526 48244 53564
rect 48860 52948 48916 53678
rect 48860 52882 48916 52892
rect 49308 54290 49924 54292
rect 49308 54238 49870 54290
rect 49922 54238 49924 54290
rect 49308 54236 49924 54238
rect 49308 52050 49364 54236
rect 49868 54226 49924 54236
rect 49532 53620 49588 53630
rect 49532 53526 49588 53564
rect 50876 53508 50932 54574
rect 50988 54516 51044 54526
rect 50988 54422 51044 54460
rect 52108 54514 52164 54908
rect 52108 54462 52110 54514
rect 52162 54462 52164 54514
rect 52108 54450 52164 54462
rect 51772 54292 51828 54302
rect 51772 54198 51828 54236
rect 52220 53956 52276 56252
rect 52108 53900 52276 53956
rect 51660 53842 51716 53854
rect 51660 53790 51662 53842
rect 51714 53790 51716 53842
rect 51660 53732 51716 53790
rect 51660 53666 51716 53676
rect 52108 53730 52164 53900
rect 52332 53844 52388 61292
rect 52444 60676 52500 60686
rect 52444 59106 52500 60620
rect 52780 60004 52836 60014
rect 52780 59910 52836 59948
rect 52444 59054 52446 59106
rect 52498 59054 52500 59106
rect 52444 58996 52500 59054
rect 52444 58930 52500 58940
rect 53004 59106 53060 59118
rect 53004 59054 53006 59106
rect 53058 59054 53060 59106
rect 52668 58212 52724 58222
rect 53004 58212 53060 59054
rect 52668 58210 53060 58212
rect 52668 58158 52670 58210
rect 52722 58158 53060 58210
rect 52668 58156 53060 58158
rect 52668 56642 52724 58156
rect 53116 57762 53172 57774
rect 53116 57710 53118 57762
rect 53170 57710 53172 57762
rect 53004 57652 53060 57662
rect 53004 57558 53060 57596
rect 52668 56590 52670 56642
rect 52722 56590 52724 56642
rect 52668 56308 52724 56590
rect 52668 56242 52724 56252
rect 52780 57540 52836 57550
rect 52108 53678 52110 53730
rect 52162 53678 52164 53730
rect 50876 53442 50932 53452
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 52108 53172 52164 53678
rect 52108 53106 52164 53116
rect 52220 53788 52388 53844
rect 52444 55188 52500 55198
rect 52556 55188 52612 55198
rect 52500 55186 52612 55188
rect 52500 55134 52558 55186
rect 52610 55134 52612 55186
rect 52500 55132 52612 55134
rect 49532 52948 49588 52958
rect 49532 52854 49588 52892
rect 50316 52836 50372 52846
rect 49308 51998 49310 52050
rect 49362 51998 49364 52050
rect 49308 51986 49364 51998
rect 49644 52834 50372 52836
rect 49644 52782 50318 52834
rect 50370 52782 50372 52834
rect 49644 52780 50372 52782
rect 49644 52050 49700 52780
rect 50316 52770 50372 52780
rect 49644 51998 49646 52050
rect 49698 51998 49700 52050
rect 49644 51986 49700 51998
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50988 50596 51044 50606
rect 48076 49970 48132 49980
rect 50428 50484 50484 50494
rect 49868 49476 49924 49486
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 49868 49026 49924 49420
rect 50428 49140 50484 50428
rect 50988 50482 51044 50540
rect 51548 50596 51604 50606
rect 51548 50502 51604 50540
rect 50988 50430 50990 50482
rect 51042 50430 51044 50482
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50540 49140 50596 49150
rect 50428 49138 50596 49140
rect 50428 49086 50542 49138
rect 50594 49086 50596 49138
rect 50428 49084 50596 49086
rect 50540 49074 50596 49084
rect 49868 48974 49870 49026
rect 49922 48974 49924 49026
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 49868 48244 49924 48974
rect 50428 48804 50484 48814
rect 50428 48356 50484 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50540 48356 50596 48366
rect 50428 48354 50596 48356
rect 50428 48302 50542 48354
rect 50594 48302 50596 48354
rect 50428 48300 50596 48302
rect 50540 48290 50596 48300
rect 49420 48242 49924 48244
rect 49420 48190 49870 48242
rect 49922 48190 49924 48242
rect 49420 48188 49924 48190
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 49420 47458 49476 48188
rect 49868 48178 49924 48188
rect 50092 47572 50148 47582
rect 50092 47478 50148 47516
rect 49420 47406 49422 47458
rect 49474 47406 49476 47458
rect 49420 47394 49476 47406
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 50876 45666 50932 45678
rect 50876 45614 50878 45666
rect 50930 45614 50932 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50764 45220 50820 45230
rect 50876 45220 50932 45614
rect 50764 45218 50932 45220
rect 50764 45166 50766 45218
rect 50818 45166 50932 45218
rect 50764 45164 50932 45166
rect 50764 45154 50820 45164
rect 50092 45106 50148 45118
rect 50092 45054 50094 45106
rect 50146 45054 50148 45106
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 49084 44322 49140 44334
rect 49084 44270 49086 44322
rect 49138 44270 49140 44322
rect 48748 44212 48804 44222
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 48748 43762 48804 44156
rect 49084 44100 49140 44270
rect 49756 44212 49812 44222
rect 49756 44118 49812 44156
rect 49084 44034 49140 44044
rect 50092 44100 50148 45054
rect 48748 43710 48750 43762
rect 48802 43710 48804 43762
rect 48748 43698 48804 43710
rect 50092 43708 50148 44044
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 49980 43652 50148 43708
rect 50988 43708 51044 50430
rect 51884 50372 51940 50382
rect 51884 50278 51940 50316
rect 51884 49810 51940 49822
rect 51884 49758 51886 49810
rect 51938 49758 51940 49810
rect 51884 49476 51940 49758
rect 51884 49410 51940 49420
rect 52220 49140 52276 53788
rect 52444 53620 52500 55132
rect 52556 55122 52612 55132
rect 52780 54516 52836 57484
rect 53116 55524 53172 57710
rect 53116 55458 53172 55468
rect 52892 54628 52948 54638
rect 52892 54626 53060 54628
rect 52892 54574 52894 54626
rect 52946 54574 53060 54626
rect 52892 54572 53060 54574
rect 52892 54562 52948 54572
rect 52780 54068 52836 54460
rect 52780 54002 52836 54012
rect 52332 53564 52500 53620
rect 53004 53732 53060 54572
rect 52332 50708 52388 53564
rect 52556 53508 52612 53518
rect 52444 52836 52500 52846
rect 52556 52836 52612 53452
rect 52892 53172 52948 53182
rect 52892 53078 52948 53116
rect 53004 52948 53060 53676
rect 53004 52882 53060 52892
rect 53116 54516 53172 54526
rect 52444 52834 52612 52836
rect 52444 52782 52446 52834
rect 52498 52782 52612 52834
rect 52444 52780 52612 52782
rect 52444 52770 52500 52780
rect 52556 52164 52612 52780
rect 52556 52098 52612 52108
rect 52892 52276 52948 52286
rect 52332 50642 52388 50652
rect 52332 50484 52388 50494
rect 52332 50390 52388 50428
rect 52668 50482 52724 50494
rect 52668 50430 52670 50482
rect 52722 50430 52724 50482
rect 52556 50372 52612 50382
rect 52108 49084 52276 49140
rect 52444 50370 52612 50372
rect 52444 50318 52558 50370
rect 52610 50318 52612 50370
rect 52444 50316 52612 50318
rect 51212 45778 51268 45790
rect 51212 45726 51214 45778
rect 51266 45726 51268 45778
rect 51212 43708 51268 45726
rect 51884 44434 51940 44446
rect 51884 44382 51886 44434
rect 51938 44382 51940 44434
rect 51884 43708 51940 44382
rect 48524 43540 48580 43550
rect 48524 43446 48580 43484
rect 49756 43540 49812 43550
rect 49756 43446 49812 43484
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 49756 42756 49812 42766
rect 49980 42756 50036 43652
rect 50764 43650 50820 43662
rect 50988 43652 51156 43708
rect 51212 43652 51716 43708
rect 51884 43652 52052 43708
rect 50764 43598 50766 43650
rect 50818 43598 50820 43650
rect 50092 43428 50148 43438
rect 50092 43334 50148 43372
rect 50764 43316 50820 43598
rect 50876 43540 50932 43550
rect 50876 43446 50932 43484
rect 50764 43250 50820 43260
rect 49756 42754 50036 42756
rect 49756 42702 49758 42754
rect 49810 42702 50036 42754
rect 49756 42700 50036 42702
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 49644 41972 49700 41982
rect 49756 41972 49812 42700
rect 50540 42644 50596 42654
rect 49644 41970 49812 41972
rect 49644 41918 49646 41970
rect 49698 41918 49812 41970
rect 49644 41916 49812 41918
rect 50428 42642 50596 42644
rect 50428 42590 50542 42642
rect 50594 42590 50596 42642
rect 50428 42588 50596 42590
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 49532 41076 49588 41086
rect 49532 40982 49588 41020
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 14252 39396 14308 39406
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2156 37886 2158 37938
rect 2210 37886 2212 37938
rect 2156 37874 2212 37886
rect 1820 37398 1876 37436
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 1820 12850 1876 12862
rect 1820 12798 1822 12850
rect 1874 12798 1876 12850
rect 1820 12516 1876 12798
rect 2156 12740 2212 12750
rect 2156 12646 2212 12684
rect 1820 12402 1876 12460
rect 1820 12350 1822 12402
rect 1874 12350 1876 12402
rect 1820 12338 1876 12350
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 6188 3444 6244 3454
rect 6636 3444 6692 3454
rect 6188 3442 6692 3444
rect 6188 3390 6190 3442
rect 6242 3390 6638 3442
rect 6690 3390 6692 3442
rect 6188 3388 6692 3390
rect 6188 3378 6244 3388
rect 6412 800 6468 3388
rect 6636 3378 6692 3388
rect 6972 3332 7028 3342
rect 6972 3238 7028 3276
rect 14252 3332 14308 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 48972 38050 49028 38062
rect 48972 37998 48974 38050
rect 49026 37998 49028 38050
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 48972 36708 49028 37998
rect 49644 38052 49700 41916
rect 50316 41860 50372 41870
rect 49868 41858 50372 41860
rect 49868 41806 50318 41858
rect 50370 41806 50372 41858
rect 49868 41804 50372 41806
rect 49868 41074 49924 41804
rect 50316 41794 50372 41804
rect 49868 41022 49870 41074
rect 49922 41022 49924 41074
rect 49868 41010 49924 41022
rect 50428 41074 50484 42588
rect 50540 42578 50596 42588
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50764 41188 50820 41198
rect 50764 41094 50820 41132
rect 50428 41022 50430 41074
rect 50482 41022 50484 41074
rect 50428 41010 50484 41022
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 51100 39506 51156 43652
rect 51660 43650 51716 43652
rect 51660 43598 51662 43650
rect 51714 43598 51716 43650
rect 51660 43586 51716 43598
rect 51996 43428 52052 43652
rect 51996 43334 52052 43372
rect 51772 41860 51828 41870
rect 51772 41410 51828 41804
rect 51772 41358 51774 41410
rect 51826 41358 51828 41410
rect 51772 41346 51828 41358
rect 51436 41076 51492 41086
rect 51436 40982 51492 41020
rect 51100 39454 51102 39506
rect 51154 39454 51156 39506
rect 50540 39396 50596 39434
rect 50540 39330 50596 39340
rect 51100 39396 51156 39454
rect 51436 39508 51492 39518
rect 51436 39414 51492 39452
rect 51100 39330 51156 39340
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50316 38946 50372 38958
rect 50316 38894 50318 38946
rect 50370 38894 50372 38946
rect 50316 38164 50372 38894
rect 52108 38948 52164 49084
rect 52444 48468 52500 50316
rect 52556 50306 52612 50316
rect 52668 49924 52724 50430
rect 52668 49858 52724 49868
rect 52556 49700 52612 49710
rect 52556 49698 52836 49700
rect 52556 49646 52558 49698
rect 52610 49646 52836 49698
rect 52556 49644 52836 49646
rect 52556 49634 52612 49644
rect 52444 48402 52500 48412
rect 52556 49476 52612 49486
rect 52220 48356 52276 48366
rect 52220 47570 52276 48300
rect 52220 47518 52222 47570
rect 52274 47518 52276 47570
rect 52220 47506 52276 47518
rect 52556 47236 52612 49420
rect 52668 49140 52724 49150
rect 52668 49046 52724 49084
rect 52780 48580 52836 49644
rect 52780 48514 52836 48524
rect 52668 48132 52724 48142
rect 52668 48038 52724 48076
rect 52668 47236 52724 47246
rect 52556 47234 52724 47236
rect 52556 47182 52670 47234
rect 52722 47182 52724 47234
rect 52556 47180 52724 47182
rect 52444 46564 52500 46574
rect 52668 46564 52724 47180
rect 52892 46788 52948 52220
rect 53116 51604 53172 54460
rect 53004 51602 53172 51604
rect 53004 51550 53118 51602
rect 53170 51550 53172 51602
rect 53004 51548 53172 51550
rect 53004 50372 53060 51548
rect 53116 51538 53172 51548
rect 53228 50484 53284 62132
rect 53340 61348 53396 61358
rect 53676 61348 53732 62974
rect 54124 62692 54180 63084
rect 54460 63140 54516 63150
rect 54460 63046 54516 63084
rect 54684 63026 54740 64540
rect 54684 62974 54686 63026
rect 54738 62974 54740 63026
rect 54684 62962 54740 62974
rect 54124 62626 54180 62636
rect 53396 61292 53732 61348
rect 53340 61254 53396 61292
rect 54908 60900 54964 67564
rect 55244 66388 55300 66398
rect 55244 65714 55300 66332
rect 55244 65662 55246 65714
rect 55298 65662 55300 65714
rect 55244 65650 55300 65662
rect 55020 65604 55076 65614
rect 55020 65510 55076 65548
rect 55356 65492 55412 65502
rect 55412 65436 55524 65492
rect 55356 65398 55412 65436
rect 55468 64818 55524 65436
rect 55468 64766 55470 64818
rect 55522 64766 55524 64818
rect 55468 64754 55524 64766
rect 55020 64482 55076 64494
rect 55020 64430 55022 64482
rect 55074 64430 55076 64482
rect 55020 63924 55076 64430
rect 55356 64372 55412 64382
rect 55020 63858 55076 63868
rect 55132 63924 55188 63934
rect 55356 63924 55412 64316
rect 55132 63922 55412 63924
rect 55132 63870 55134 63922
rect 55186 63870 55412 63922
rect 55132 63868 55412 63870
rect 55132 63858 55188 63868
rect 55356 63138 55412 63868
rect 55356 63086 55358 63138
rect 55410 63086 55412 63138
rect 55356 63074 55412 63086
rect 55132 62580 55188 62590
rect 55132 61794 55188 62524
rect 55356 62356 55412 62366
rect 55580 62356 55636 70140
rect 55692 69524 55748 69534
rect 55692 63922 55748 69468
rect 56252 68626 56308 70364
rect 56476 70306 56532 70476
rect 56476 70254 56478 70306
rect 56530 70254 56532 70306
rect 56476 70242 56532 70254
rect 56476 69524 56532 69534
rect 56476 69430 56532 69468
rect 57148 69524 57204 69534
rect 57148 69410 57204 69468
rect 57148 69358 57150 69410
rect 57202 69358 57204 69410
rect 57148 69346 57204 69358
rect 56476 69300 56532 69310
rect 56476 68850 56532 69244
rect 57372 68852 57428 70588
rect 57596 69972 57652 69982
rect 57596 69878 57652 69916
rect 57932 69970 57988 69982
rect 57932 69918 57934 69970
rect 57986 69918 57988 69970
rect 57932 69636 57988 69918
rect 57932 69570 57988 69580
rect 57820 69300 57876 69310
rect 57820 69206 57876 69244
rect 56476 68798 56478 68850
rect 56530 68798 56532 68850
rect 56476 68786 56532 68798
rect 57036 68850 57428 68852
rect 57036 68798 57374 68850
rect 57426 68798 57428 68850
rect 57036 68796 57428 68798
rect 56252 68574 56254 68626
rect 56306 68574 56308 68626
rect 56252 68562 56308 68574
rect 56476 66388 56532 66398
rect 56476 66294 56532 66332
rect 57036 66386 57092 68796
rect 57372 68786 57428 68796
rect 57036 66334 57038 66386
rect 57090 66334 57092 66386
rect 57036 66322 57092 66334
rect 58044 66388 58100 66398
rect 55804 66276 55860 66286
rect 55804 65492 55860 66220
rect 55804 65360 55860 65436
rect 57596 65490 57652 65502
rect 57596 65438 57598 65490
rect 57650 65438 57652 65490
rect 56700 65378 56756 65390
rect 56700 65326 56702 65378
rect 56754 65326 56756 65378
rect 56364 64820 56420 64830
rect 56700 64820 56756 65326
rect 56700 64764 57092 64820
rect 56364 64726 56420 64764
rect 56924 64594 56980 64606
rect 56924 64542 56926 64594
rect 56978 64542 56980 64594
rect 55692 63870 55694 63922
rect 55746 63870 55748 63922
rect 55692 63858 55748 63870
rect 56364 64482 56420 64494
rect 56364 64430 56366 64482
rect 56418 64430 56420 64482
rect 55692 63476 55748 63486
rect 55692 63138 55748 63420
rect 56364 63476 56420 64430
rect 56476 64484 56532 64494
rect 56476 64390 56532 64428
rect 56700 64482 56756 64494
rect 56700 64430 56702 64482
rect 56754 64430 56756 64482
rect 56700 64036 56756 64430
rect 56924 64260 56980 64542
rect 56924 64194 56980 64204
rect 56700 63980 56980 64036
rect 56588 63924 56644 63934
rect 56588 63922 56868 63924
rect 56588 63870 56590 63922
rect 56642 63870 56868 63922
rect 56588 63868 56868 63870
rect 56588 63858 56644 63868
rect 56364 63410 56420 63420
rect 56700 63140 56756 63150
rect 55692 63086 55694 63138
rect 55746 63086 55748 63138
rect 55692 63074 55748 63086
rect 56252 63138 56756 63140
rect 56252 63086 56702 63138
rect 56754 63086 56756 63138
rect 56252 63084 56756 63086
rect 55804 62356 55860 62366
rect 55356 62354 55860 62356
rect 55356 62302 55358 62354
rect 55410 62302 55806 62354
rect 55858 62302 55860 62354
rect 55356 62300 55860 62302
rect 55356 62290 55412 62300
rect 55804 62290 55860 62300
rect 55132 61742 55134 61794
rect 55186 61742 55188 61794
rect 55132 61730 55188 61742
rect 56140 61572 56196 61582
rect 55020 61460 55076 61470
rect 55020 61366 55076 61404
rect 55692 61460 55748 61470
rect 55692 61366 55748 61404
rect 55132 61348 55188 61358
rect 55132 61254 55188 61292
rect 56140 61348 56196 61516
rect 56140 61254 56196 61292
rect 56252 61012 56308 63084
rect 56700 63074 56756 63084
rect 56700 62692 56756 62702
rect 56700 62578 56756 62636
rect 56700 62526 56702 62578
rect 56754 62526 56756 62578
rect 56700 62514 56756 62526
rect 56252 61010 56644 61012
rect 56252 60958 56254 61010
rect 56306 60958 56644 61010
rect 56252 60956 56644 60958
rect 56252 60946 56308 60956
rect 54236 60844 54964 60900
rect 55468 60898 55524 60910
rect 55468 60846 55470 60898
rect 55522 60846 55524 60898
rect 53676 60004 53732 60014
rect 53676 59910 53732 59948
rect 53788 59218 53844 59230
rect 53788 59166 53790 59218
rect 53842 59166 53844 59218
rect 53452 58210 53508 58222
rect 53452 58158 53454 58210
rect 53506 58158 53508 58210
rect 53340 57650 53396 57662
rect 53340 57598 53342 57650
rect 53394 57598 53396 57650
rect 53340 56980 53396 57598
rect 53452 57652 53508 58158
rect 53788 57652 53844 59166
rect 53452 57650 53844 57652
rect 53452 57598 53790 57650
rect 53842 57598 53844 57650
rect 53452 57596 53844 57598
rect 53340 56914 53396 56924
rect 53564 56866 53620 56878
rect 53564 56814 53566 56866
rect 53618 56814 53620 56866
rect 53564 56308 53620 56814
rect 53788 56308 53844 57596
rect 53620 56252 53844 56308
rect 53564 56242 53620 56252
rect 53788 55298 53844 56252
rect 54236 59220 54292 60844
rect 55244 60788 55300 60798
rect 54572 60786 55300 60788
rect 54572 60734 55246 60786
rect 55298 60734 55300 60786
rect 54572 60732 55300 60734
rect 54460 59890 54516 59902
rect 54460 59838 54462 59890
rect 54514 59838 54516 59890
rect 54236 55468 54292 59164
rect 54348 59668 54404 59678
rect 54348 58434 54404 59612
rect 54460 59444 54516 59838
rect 54460 59378 54516 59388
rect 54572 59330 54628 60732
rect 55244 60722 55300 60732
rect 54572 59278 54574 59330
rect 54626 59278 54628 59330
rect 54572 59266 54628 59278
rect 55468 58884 55524 60846
rect 55580 60786 55636 60798
rect 55580 60734 55582 60786
rect 55634 60734 55636 60786
rect 55580 60228 55636 60734
rect 56140 60788 56196 60798
rect 56140 60694 56196 60732
rect 56476 60786 56532 60798
rect 56476 60734 56478 60786
rect 56530 60734 56532 60786
rect 55580 60162 55636 60172
rect 56476 59556 56532 60734
rect 56588 60114 56644 60956
rect 56588 60062 56590 60114
rect 56642 60062 56644 60114
rect 56588 60050 56644 60062
rect 56812 59892 56868 63868
rect 56924 63140 56980 63980
rect 56924 63074 56980 63084
rect 57036 62692 57092 64764
rect 57596 64708 57652 65438
rect 57596 64642 57652 64652
rect 57820 65490 57876 65502
rect 57820 65438 57822 65490
rect 57874 65438 57876 65490
rect 57484 64596 57540 64606
rect 57484 64502 57540 64540
rect 57820 64596 57876 65438
rect 57708 64482 57764 64494
rect 57708 64430 57710 64482
rect 57762 64430 57764 64482
rect 57596 64372 57652 64382
rect 57484 64036 57540 64046
rect 57484 63942 57540 63980
rect 57596 63812 57652 64316
rect 57484 63756 57652 63812
rect 57036 62626 57092 62636
rect 57372 63364 57428 63374
rect 57372 62354 57428 63308
rect 57484 63250 57540 63756
rect 57484 63198 57486 63250
rect 57538 63198 57540 63250
rect 57484 63186 57540 63198
rect 57596 63476 57652 63486
rect 57596 62578 57652 63420
rect 57708 63364 57764 64430
rect 57708 63298 57764 63308
rect 57596 62526 57598 62578
rect 57650 62526 57652 62578
rect 57596 62514 57652 62526
rect 57372 62302 57374 62354
rect 57426 62302 57428 62354
rect 57372 62290 57428 62302
rect 57820 62466 57876 64540
rect 57932 65378 57988 65390
rect 57932 65326 57934 65378
rect 57986 65326 57988 65378
rect 57932 64148 57988 65326
rect 58044 65268 58100 66332
rect 58268 66388 58324 71820
rect 58492 71652 58548 71662
rect 58492 70306 58548 71596
rect 58828 71650 58884 71662
rect 58828 71598 58830 71650
rect 58882 71598 58884 71650
rect 58604 70754 58660 70766
rect 58604 70702 58606 70754
rect 58658 70702 58660 70754
rect 58604 70420 58660 70702
rect 58604 70354 58660 70364
rect 58492 70254 58494 70306
rect 58546 70254 58548 70306
rect 58492 70242 58548 70254
rect 58716 70194 58772 70206
rect 58716 70142 58718 70194
rect 58770 70142 58772 70194
rect 58716 70084 58772 70142
rect 58828 70196 58884 71598
rect 59052 71092 59108 72382
rect 59052 71026 59108 71036
rect 58828 70130 58884 70140
rect 58940 70978 58996 70990
rect 58940 70926 58942 70978
rect 58994 70926 58996 70978
rect 58716 68852 58772 70028
rect 58940 69972 58996 70926
rect 59164 70866 59220 72494
rect 59164 70814 59166 70866
rect 59218 70814 59220 70866
rect 59164 70802 59220 70814
rect 59500 71092 59556 71102
rect 59500 70866 59556 71036
rect 59500 70814 59502 70866
rect 59554 70814 59556 70866
rect 59500 70802 59556 70814
rect 59836 70308 59892 73892
rect 60396 72548 60452 72558
rect 60396 72454 60452 72492
rect 60284 70754 60340 70766
rect 60284 70702 60286 70754
rect 60338 70702 60340 70754
rect 60284 70644 60340 70702
rect 60508 70644 60564 78932
rect 61292 78596 61348 78606
rect 61292 78502 61348 78540
rect 60956 78372 61012 78382
rect 60956 78034 61012 78316
rect 60956 77982 60958 78034
rect 61010 77982 61012 78034
rect 60956 77970 61012 77982
rect 61516 78034 61572 80556
rect 61628 79490 61684 79502
rect 61628 79438 61630 79490
rect 61682 79438 61684 79490
rect 61628 78988 61684 79438
rect 61628 78932 61796 78988
rect 61740 78594 61796 78932
rect 61740 78542 61742 78594
rect 61794 78542 61796 78594
rect 61740 78372 61796 78542
rect 61740 78306 61796 78316
rect 61516 77982 61518 78034
rect 61570 77982 61572 78034
rect 61516 77970 61572 77982
rect 62188 78036 62244 81900
rect 62412 78988 62468 85708
rect 62972 86658 63028 86670
rect 62972 86606 62974 86658
rect 63026 86606 63028 86658
rect 62972 85764 63028 86606
rect 63420 86212 63476 87166
rect 63420 86146 63476 86156
rect 63084 85876 63140 85886
rect 63084 85782 63140 85820
rect 62972 85698 63028 85708
rect 62636 85204 62692 85214
rect 62524 85202 62692 85204
rect 62524 85150 62638 85202
rect 62690 85150 62692 85202
rect 62524 85148 62692 85150
rect 62524 81956 62580 85148
rect 62636 85138 62692 85148
rect 63420 83748 63476 83758
rect 63532 83748 63588 88062
rect 63868 88004 63924 88014
rect 63868 88002 64260 88004
rect 63868 87950 63870 88002
rect 63922 87950 64260 88002
rect 63868 87948 64260 87950
rect 63868 87938 63924 87948
rect 63756 87220 63812 87230
rect 63756 87126 63812 87164
rect 63420 83746 63588 83748
rect 63420 83694 63422 83746
rect 63474 83694 63588 83746
rect 63420 83692 63588 83694
rect 63644 86546 63700 86558
rect 63644 86494 63646 86546
rect 63698 86494 63700 86546
rect 63420 83682 63476 83692
rect 63644 83524 63700 86494
rect 64204 86548 64260 87948
rect 64428 88002 64484 88014
rect 64428 87950 64430 88002
rect 64482 87950 64484 88002
rect 64428 87892 64484 87950
rect 64428 87826 64484 87836
rect 64316 87556 64372 87566
rect 64316 87462 64372 87500
rect 64540 87444 64596 87454
rect 65324 87444 65380 87454
rect 64540 87442 65380 87444
rect 64540 87390 64542 87442
rect 64594 87390 65326 87442
rect 65378 87390 65380 87442
rect 64540 87388 65380 87390
rect 64540 87378 64596 87388
rect 64204 86492 64820 86548
rect 64540 86324 64596 86334
rect 63868 85874 63924 85886
rect 63868 85822 63870 85874
rect 63922 85822 63924 85874
rect 63868 85764 63924 85822
rect 63868 85698 63924 85708
rect 64316 85764 64372 85774
rect 64316 85670 64372 85708
rect 63756 84868 63812 84878
rect 63756 83748 63812 84812
rect 64316 84308 64372 84318
rect 64316 84214 64372 84252
rect 64428 84084 64484 84094
rect 63756 83692 63924 83748
rect 63420 83468 63700 83524
rect 63756 83522 63812 83534
rect 63756 83470 63758 83522
rect 63810 83470 63812 83522
rect 63420 82962 63476 83468
rect 63756 83412 63812 83470
rect 63420 82910 63422 82962
rect 63474 82910 63476 82962
rect 63420 82898 63476 82910
rect 63644 83356 63812 83412
rect 62524 81890 62580 81900
rect 62636 81954 62692 81966
rect 62636 81902 62638 81954
rect 62690 81902 62692 81954
rect 62636 80612 62692 81902
rect 63420 81954 63476 81966
rect 63420 81902 63422 81954
rect 63474 81902 63476 81954
rect 63196 81844 63252 81854
rect 62636 80546 62692 80556
rect 62972 81842 63252 81844
rect 62972 81790 63198 81842
rect 63250 81790 63252 81842
rect 62972 81788 63252 81790
rect 62972 80500 63028 81788
rect 63196 81778 63252 81788
rect 63420 81732 63476 81902
rect 63644 81956 63700 83356
rect 63868 83300 63924 83692
rect 64428 83522 64484 84028
rect 64428 83470 64430 83522
rect 64482 83470 64484 83522
rect 64428 83458 64484 83470
rect 64540 83410 64596 86268
rect 64764 85202 64820 86492
rect 64764 85150 64766 85202
rect 64818 85150 64820 85202
rect 64764 85138 64820 85150
rect 65100 84084 65156 87388
rect 65324 87378 65380 87388
rect 67452 87442 67508 87454
rect 67452 87390 67454 87442
rect 67506 87390 67508 87442
rect 67452 87332 67508 87390
rect 65916 87052 66180 87062
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 65916 86986 66180 86996
rect 65772 86770 65828 86782
rect 65772 86718 65774 86770
rect 65826 86718 65828 86770
rect 65548 86436 65604 86446
rect 65436 85764 65492 85774
rect 65548 85764 65604 86380
rect 65772 86324 65828 86718
rect 65772 85876 65828 86268
rect 66332 86434 66388 86446
rect 66332 86382 66334 86434
rect 66386 86382 66388 86434
rect 66332 85876 66388 86382
rect 66668 86436 66724 86446
rect 66668 86342 66724 86380
rect 66444 85876 66500 85886
rect 66332 85874 66500 85876
rect 66332 85822 66446 85874
rect 66498 85822 66500 85874
rect 66332 85820 66500 85822
rect 65772 85810 65828 85820
rect 65492 85708 65604 85764
rect 65436 85632 65492 85708
rect 65548 85092 65604 85708
rect 65916 85484 66180 85494
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 65916 85418 66180 85428
rect 65548 85090 65940 85092
rect 65548 85038 65550 85090
rect 65602 85038 65940 85090
rect 65548 85036 65940 85038
rect 65548 85026 65604 85036
rect 65772 84532 65828 84542
rect 65100 83634 65156 84028
rect 65100 83582 65102 83634
rect 65154 83582 65156 83634
rect 65100 83570 65156 83582
rect 65660 84476 65772 84532
rect 64540 83358 64542 83410
rect 64594 83358 64596 83410
rect 64540 83346 64596 83358
rect 63756 83244 63924 83300
rect 63756 82850 63812 83244
rect 63756 82798 63758 82850
rect 63810 82798 63812 82850
rect 63756 82786 63812 82798
rect 63980 82068 64036 82078
rect 63980 81974 64036 82012
rect 63644 81890 63700 81900
rect 62748 79716 62804 79726
rect 62972 79716 63028 80444
rect 63308 81676 63420 81732
rect 63308 80164 63364 81676
rect 63420 81666 63476 81676
rect 64092 81732 64148 81742
rect 63980 81284 64036 81294
rect 63532 81282 64036 81284
rect 63532 81230 63982 81282
rect 64034 81230 64036 81282
rect 63532 81228 64036 81230
rect 63420 81058 63476 81070
rect 63420 81006 63422 81058
rect 63474 81006 63476 81058
rect 63420 80612 63476 81006
rect 63420 80546 63476 80556
rect 63532 80498 63588 81228
rect 63980 81218 64036 81228
rect 63532 80446 63534 80498
rect 63586 80446 63588 80498
rect 63532 80434 63588 80446
rect 63644 80724 63700 80734
rect 62748 79714 63028 79716
rect 62748 79662 62750 79714
rect 62802 79662 63028 79714
rect 62748 79660 63028 79662
rect 63084 80108 63364 80164
rect 63084 79714 63140 80108
rect 63644 79826 63700 80668
rect 64092 80164 64148 81676
rect 64428 81732 64484 81742
rect 64428 81638 64484 81676
rect 64204 81170 64260 81182
rect 64204 81118 64206 81170
rect 64258 81118 64260 81170
rect 64204 80724 64260 81118
rect 64204 80658 64260 80668
rect 64316 80388 64372 80398
rect 64316 80386 64484 80388
rect 64316 80334 64318 80386
rect 64370 80334 64484 80386
rect 64316 80332 64484 80334
rect 64316 80322 64372 80332
rect 64428 80164 64484 80332
rect 64764 80164 64820 80174
rect 64092 80108 64372 80164
rect 63644 79774 63646 79826
rect 63698 79774 63700 79826
rect 63644 79762 63700 79774
rect 64316 79826 64372 80108
rect 64316 79774 64318 79826
rect 64370 79774 64372 79826
rect 64316 79762 64372 79774
rect 64428 80162 64820 80164
rect 64428 80110 64766 80162
rect 64818 80110 64820 80162
rect 64428 80108 64820 80110
rect 63084 79662 63086 79714
rect 63138 79662 63140 79714
rect 62748 79650 62804 79660
rect 63084 79650 63140 79662
rect 62300 78932 62468 78988
rect 62636 79604 62692 79614
rect 62300 78820 62356 78932
rect 62300 78726 62356 78764
rect 62636 78594 62692 79548
rect 63308 79604 63364 79614
rect 63308 79510 63364 79548
rect 64316 78820 64372 78830
rect 63980 78818 64372 78820
rect 63980 78766 64318 78818
rect 64370 78766 64372 78818
rect 63980 78764 64372 78766
rect 62636 78542 62638 78594
rect 62690 78542 62692 78594
rect 62300 78036 62356 78046
rect 62188 78034 62356 78036
rect 62188 77982 62302 78034
rect 62354 77982 62356 78034
rect 62188 77980 62356 77982
rect 62300 77970 62356 77980
rect 61628 77700 61684 77710
rect 61516 75908 61572 75918
rect 60620 74900 60676 74910
rect 60620 74806 60676 74844
rect 61292 74788 61348 74798
rect 60732 74786 61348 74788
rect 60732 74734 61294 74786
rect 61346 74734 61348 74786
rect 60732 74732 61348 74734
rect 60620 74004 60676 74014
rect 60732 74004 60788 74732
rect 61292 74722 61348 74732
rect 61516 74788 61572 75852
rect 61516 74722 61572 74732
rect 61516 74116 61572 74126
rect 61516 74022 61572 74060
rect 60620 74002 60788 74004
rect 60620 73950 60622 74002
rect 60674 73950 60788 74002
rect 60620 73948 60788 73950
rect 60620 73938 60676 73948
rect 61516 73556 61572 73566
rect 61516 73330 61572 73500
rect 61516 73278 61518 73330
rect 61570 73278 61572 73330
rect 61516 73266 61572 73278
rect 60844 73220 60900 73230
rect 60844 73126 60900 73164
rect 60620 72322 60676 72334
rect 60620 72270 60622 72322
rect 60674 72270 60676 72322
rect 60620 71092 60676 72270
rect 60620 71026 60676 71036
rect 60956 71204 61012 71214
rect 60508 70588 60900 70644
rect 60284 70578 60340 70588
rect 59388 70252 59892 70308
rect 60620 70420 60676 70430
rect 59276 70196 59332 70206
rect 59276 70102 59332 70140
rect 59052 69972 59108 69982
rect 58940 69970 59108 69972
rect 58940 69918 59054 69970
rect 59106 69918 59108 69970
rect 58940 69916 59108 69918
rect 59052 69906 59108 69916
rect 58716 68786 58772 68796
rect 59388 67956 59444 70252
rect 60620 70196 60676 70364
rect 60396 70194 60676 70196
rect 60396 70142 60622 70194
rect 60674 70142 60676 70194
rect 60396 70140 60676 70142
rect 59724 70084 59780 70094
rect 59724 69990 59780 70028
rect 59836 69970 59892 69982
rect 59836 69918 59838 69970
rect 59890 69918 59892 69970
rect 59836 69748 59892 69918
rect 58940 67954 59444 67956
rect 58940 67902 59390 67954
rect 59442 67902 59444 67954
rect 58940 67900 59444 67902
rect 58716 66948 58772 66958
rect 58716 66946 58884 66948
rect 58716 66894 58718 66946
rect 58770 66894 58884 66946
rect 58716 66892 58884 66894
rect 58716 66882 58772 66892
rect 58268 66386 58772 66388
rect 58268 66334 58270 66386
rect 58322 66334 58772 66386
rect 58268 66332 58772 66334
rect 58268 66322 58324 66332
rect 58604 66052 58660 66062
rect 58492 66050 58660 66052
rect 58492 65998 58606 66050
rect 58658 65998 58660 66050
rect 58492 65996 58660 65998
rect 58156 65492 58212 65502
rect 58156 65490 58436 65492
rect 58156 65438 58158 65490
rect 58210 65438 58436 65490
rect 58156 65436 58436 65438
rect 58156 65426 58212 65436
rect 58044 65212 58212 65268
rect 57932 64082 57988 64092
rect 58044 64708 58100 64718
rect 57932 63924 57988 63934
rect 57932 63830 57988 63868
rect 58044 63700 58100 64652
rect 58156 63924 58212 65212
rect 58380 64148 58436 65436
rect 58492 64708 58548 65996
rect 58604 65986 58660 65996
rect 58716 65828 58772 66332
rect 58828 66164 58884 66892
rect 58940 66274 58996 67900
rect 59388 67890 59444 67900
rect 59724 69692 60004 69748
rect 58940 66222 58942 66274
rect 58994 66222 58996 66274
rect 58940 66210 58996 66222
rect 59052 66946 59108 66958
rect 59052 66894 59054 66946
rect 59106 66894 59108 66946
rect 58828 66032 58884 66108
rect 58604 65772 58772 65828
rect 58828 65828 58884 65838
rect 58604 65602 58660 65772
rect 58604 65550 58606 65602
rect 58658 65550 58660 65602
rect 58604 65538 58660 65550
rect 58716 65604 58772 65614
rect 58828 65604 58884 65772
rect 59052 65828 59108 66894
rect 59052 65762 59108 65772
rect 59500 66050 59556 66062
rect 59500 65998 59502 66050
rect 59554 65998 59556 66050
rect 58716 65602 58884 65604
rect 58716 65550 58718 65602
rect 58770 65550 58884 65602
rect 58716 65548 58884 65550
rect 58716 65538 58772 65548
rect 58940 65492 58996 65502
rect 58940 65398 58996 65436
rect 59276 65380 59332 65390
rect 59276 65378 59444 65380
rect 59276 65326 59278 65378
rect 59330 65326 59444 65378
rect 59276 65324 59444 65326
rect 59276 65314 59332 65324
rect 58492 64652 58660 64708
rect 58492 64482 58548 64494
rect 58492 64430 58494 64482
rect 58546 64430 58548 64482
rect 58492 64372 58548 64430
rect 58492 64306 58548 64316
rect 58492 64148 58548 64158
rect 58380 64146 58548 64148
rect 58380 64094 58494 64146
rect 58546 64094 58548 64146
rect 58380 64092 58548 64094
rect 58492 64082 58548 64092
rect 58268 63924 58324 63934
rect 58156 63922 58324 63924
rect 58156 63870 58270 63922
rect 58322 63870 58324 63922
rect 58156 63868 58324 63870
rect 58268 63858 58324 63868
rect 57820 62414 57822 62466
rect 57874 62414 57876 62466
rect 57820 62356 57876 62414
rect 57820 62290 57876 62300
rect 57932 63644 58100 63700
rect 57932 62354 57988 63644
rect 58156 63364 58212 63374
rect 58156 63138 58212 63308
rect 58268 63252 58324 63262
rect 58268 63158 58324 63196
rect 58156 63086 58158 63138
rect 58210 63086 58212 63138
rect 58156 63074 58212 63086
rect 58380 63140 58436 63150
rect 58604 63140 58660 64652
rect 59388 64596 59444 65324
rect 59500 64708 59556 65998
rect 59500 64642 59556 64652
rect 59612 65492 59668 65502
rect 59388 64502 59444 64540
rect 58940 64482 58996 64494
rect 58940 64430 58942 64482
rect 58994 64430 58996 64482
rect 58380 63138 58660 63140
rect 58380 63086 58382 63138
rect 58434 63086 58660 63138
rect 58380 63084 58660 63086
rect 58716 64036 58772 64046
rect 58380 63074 58436 63084
rect 58604 62914 58660 62926
rect 58604 62862 58606 62914
rect 58658 62862 58660 62914
rect 58604 62580 58660 62862
rect 58604 62514 58660 62524
rect 57932 62302 57934 62354
rect 57986 62302 57988 62354
rect 57932 62188 57988 62302
rect 58604 62356 58660 62366
rect 58604 62262 58660 62300
rect 57932 62132 58436 62188
rect 58380 62020 58436 62132
rect 58380 61964 58660 62020
rect 58604 61682 58660 61964
rect 58604 61630 58606 61682
rect 58658 61630 58660 61682
rect 58604 61618 58660 61630
rect 56476 59490 56532 59500
rect 56700 59836 56812 59892
rect 56700 59106 56756 59836
rect 56812 59826 56868 59836
rect 57036 61348 57092 61358
rect 56700 59054 56702 59106
rect 56754 59054 56756 59106
rect 56700 59042 56756 59054
rect 56812 59332 56868 59342
rect 55468 58818 55524 58828
rect 54348 58382 54350 58434
rect 54402 58382 54404 58434
rect 54348 58370 54404 58382
rect 54460 58660 54516 58670
rect 54460 58322 54516 58604
rect 55244 58436 55300 58446
rect 55244 58342 55300 58380
rect 54460 58270 54462 58322
rect 54514 58270 54516 58322
rect 54460 58258 54516 58270
rect 54684 58324 54740 58334
rect 54684 58230 54740 58268
rect 55916 58324 55972 58334
rect 55916 58230 55972 58268
rect 54572 57538 54628 57550
rect 54572 57486 54574 57538
rect 54626 57486 54628 57538
rect 54348 56980 54404 56990
rect 54348 56886 54404 56924
rect 54460 56420 54516 56430
rect 54236 55412 54404 55468
rect 53788 55246 53790 55298
rect 53842 55246 53844 55298
rect 53788 54740 53844 55246
rect 54348 54964 54404 55412
rect 54460 55410 54516 56364
rect 54572 56308 54628 57486
rect 56700 57540 56756 57550
rect 56812 57540 56868 59276
rect 56700 57538 56868 57540
rect 56700 57486 56702 57538
rect 56754 57486 56868 57538
rect 56700 57484 56868 57486
rect 56700 57474 56756 57484
rect 56700 57092 56756 57102
rect 56476 56978 56532 56990
rect 56476 56926 56478 56978
rect 56530 56926 56532 56978
rect 56476 56756 56532 56926
rect 56476 56690 56532 56700
rect 54572 56242 54628 56252
rect 56588 56644 56644 56654
rect 56476 56084 56532 56094
rect 56476 55990 56532 56028
rect 54460 55358 54462 55410
rect 54514 55358 54516 55410
rect 54460 55346 54516 55358
rect 55468 55524 55524 55534
rect 54348 54908 55300 54964
rect 54348 54740 54404 54750
rect 53788 54738 54404 54740
rect 53788 54686 54350 54738
rect 54402 54686 54404 54738
rect 53788 54684 54404 54686
rect 54348 54674 54404 54684
rect 55020 54516 55076 54526
rect 55020 54422 55076 54460
rect 53452 54402 53508 54414
rect 53452 54350 53454 54402
rect 53506 54350 53508 54402
rect 53452 54068 53508 54350
rect 53452 54002 53508 54012
rect 53900 54402 53956 54414
rect 53900 54350 53902 54402
rect 53954 54350 53956 54402
rect 53900 54068 53956 54350
rect 53900 54002 53956 54012
rect 55132 52948 55188 52958
rect 53340 52276 53396 52286
rect 53340 52182 53396 52220
rect 53788 52164 53844 52174
rect 54572 52164 54628 52174
rect 53788 52162 54628 52164
rect 53788 52110 53790 52162
rect 53842 52110 54574 52162
rect 54626 52110 54628 52162
rect 53788 52108 54628 52110
rect 53788 52098 53844 52108
rect 54348 51940 54404 51950
rect 54124 51716 54180 51726
rect 53676 50708 53732 50718
rect 53676 50594 53732 50652
rect 53676 50542 53678 50594
rect 53730 50542 53732 50594
rect 53676 50530 53732 50542
rect 53004 50306 53060 50316
rect 53116 50428 53284 50484
rect 53116 48468 53172 50428
rect 53340 50372 53396 50382
rect 53228 50370 53396 50372
rect 53228 50318 53342 50370
rect 53394 50318 53396 50370
rect 53228 50316 53396 50318
rect 53228 48580 53284 50316
rect 53340 50306 53396 50316
rect 53564 50372 53620 50382
rect 53564 50278 53620 50316
rect 54124 49140 54180 51660
rect 54348 51602 54404 51884
rect 54348 51550 54350 51602
rect 54402 51550 54404 51602
rect 54348 51538 54404 51550
rect 54236 51154 54292 51166
rect 54236 51102 54238 51154
rect 54290 51102 54292 51154
rect 54236 50482 54292 51102
rect 54236 50430 54238 50482
rect 54290 50430 54292 50482
rect 54236 50036 54292 50430
rect 54348 50596 54404 50606
rect 54572 50596 54628 52108
rect 55020 52162 55076 52174
rect 55020 52110 55022 52162
rect 55074 52110 55076 52162
rect 55020 51940 55076 52110
rect 55020 51874 55076 51884
rect 54796 51268 54852 51278
rect 54796 51266 54964 51268
rect 54796 51214 54798 51266
rect 54850 51214 54964 51266
rect 54796 51212 54964 51214
rect 54796 51202 54852 51212
rect 54908 50708 54964 51212
rect 54572 50540 54852 50596
rect 54348 50372 54404 50540
rect 54572 50372 54628 50382
rect 54348 50370 54516 50372
rect 54348 50318 54350 50370
rect 54402 50318 54516 50370
rect 54348 50316 54516 50318
rect 54348 50306 54404 50316
rect 54460 50148 54516 50316
rect 54572 50278 54628 50316
rect 54460 50092 54740 50148
rect 54236 49980 54516 50036
rect 54348 49812 54404 49822
rect 54348 49250 54404 49756
rect 54348 49198 54350 49250
rect 54402 49198 54404 49250
rect 54348 49186 54404 49198
rect 54460 49588 54516 49980
rect 54684 49698 54740 50092
rect 54684 49646 54686 49698
rect 54738 49646 54740 49698
rect 54684 49634 54740 49646
rect 54124 49028 54180 49084
rect 54124 48972 54404 49028
rect 53676 48914 53732 48926
rect 53676 48862 53678 48914
rect 53730 48862 53732 48914
rect 53340 48804 53396 48814
rect 53340 48710 53396 48748
rect 53564 48804 53620 48814
rect 53564 48710 53620 48748
rect 53228 48524 53396 48580
rect 53116 48412 53284 48468
rect 53116 48242 53172 48254
rect 53116 48190 53118 48242
rect 53170 48190 53172 48242
rect 53116 47572 53172 48190
rect 53116 47506 53172 47516
rect 52892 46732 53060 46788
rect 52892 46564 52948 46574
rect 52444 46562 52948 46564
rect 52444 46510 52446 46562
rect 52498 46510 52894 46562
rect 52946 46510 52948 46562
rect 52444 46508 52948 46510
rect 52444 46498 52500 46508
rect 52892 45332 52948 46508
rect 52892 45266 52948 45276
rect 52892 44996 52948 45006
rect 53004 44996 53060 46732
rect 53228 46676 53284 48412
rect 53340 48466 53396 48524
rect 53340 48414 53342 48466
rect 53394 48414 53396 48466
rect 53340 48402 53396 48414
rect 53452 48468 53508 48478
rect 53452 48354 53508 48412
rect 53452 48302 53454 48354
rect 53506 48302 53508 48354
rect 53452 48290 53508 48302
rect 53676 48244 53732 48862
rect 54348 48914 54404 48972
rect 54348 48862 54350 48914
rect 54402 48862 54404 48914
rect 54348 48850 54404 48862
rect 54460 48914 54516 49532
rect 54796 49476 54852 50540
rect 54908 50484 54964 50652
rect 55132 50596 55188 52892
rect 55244 51492 55300 54908
rect 55468 54738 55524 55468
rect 56588 55410 56644 56588
rect 56588 55358 56590 55410
rect 56642 55358 56644 55410
rect 56588 55346 56644 55358
rect 55468 54686 55470 54738
rect 55522 54686 55524 54738
rect 55468 54674 55524 54686
rect 55580 55300 55636 55310
rect 55356 52162 55412 52174
rect 55356 52110 55358 52162
rect 55410 52110 55412 52162
rect 55356 51716 55412 52110
rect 55580 52050 55636 55244
rect 56700 54738 56756 57036
rect 57036 55300 57092 61292
rect 58716 61124 58772 63980
rect 58940 64036 58996 64430
rect 59276 64372 59332 64382
rect 58940 63970 58996 63980
rect 59052 64148 59108 64158
rect 58940 63140 58996 63150
rect 59052 63140 59108 64092
rect 59164 63924 59220 63934
rect 59276 63924 59332 64316
rect 59164 63922 59332 63924
rect 59164 63870 59166 63922
rect 59218 63870 59332 63922
rect 59164 63868 59332 63870
rect 59164 63858 59220 63868
rect 59500 63588 59556 63598
rect 59500 63250 59556 63532
rect 59500 63198 59502 63250
rect 59554 63198 59556 63250
rect 59500 63186 59556 63198
rect 59388 63140 59444 63150
rect 59052 63138 59444 63140
rect 59052 63086 59390 63138
rect 59442 63086 59444 63138
rect 59052 63084 59444 63086
rect 58828 63026 58884 63038
rect 58828 62974 58830 63026
rect 58882 62974 58884 63026
rect 58828 62916 58884 62974
rect 58828 62850 58884 62860
rect 58940 61570 58996 63084
rect 59388 63074 59444 63084
rect 59612 63138 59668 65436
rect 59724 63922 59780 69692
rect 59836 69524 59892 69534
rect 59836 67060 59892 69468
rect 59948 69522 60004 69692
rect 59948 69470 59950 69522
rect 60002 69470 60004 69522
rect 59948 69458 60004 69470
rect 60396 69524 60452 70140
rect 60620 70130 60676 70140
rect 60732 70196 60788 70206
rect 60396 69392 60452 69468
rect 60732 68964 60788 70140
rect 60620 68852 60676 68862
rect 60732 68852 60788 68908
rect 60620 68850 60788 68852
rect 60620 68798 60622 68850
rect 60674 68798 60788 68850
rect 60620 68796 60788 68798
rect 60620 68786 60676 68796
rect 60620 67732 60676 67742
rect 60620 67638 60676 67676
rect 60284 67620 60340 67630
rect 60284 67618 60452 67620
rect 60284 67566 60286 67618
rect 60338 67566 60452 67618
rect 60284 67564 60452 67566
rect 60284 67554 60340 67564
rect 60396 67172 60452 67564
rect 60508 67172 60564 67182
rect 60396 67170 60564 67172
rect 60396 67118 60510 67170
rect 60562 67118 60564 67170
rect 60396 67116 60564 67118
rect 60508 67106 60564 67116
rect 59836 67058 60004 67060
rect 59836 67006 59838 67058
rect 59890 67006 60004 67058
rect 59836 67004 60004 67006
rect 59836 66994 59892 67004
rect 59948 65490 60004 67004
rect 60396 66276 60452 66286
rect 60396 66182 60452 66220
rect 59948 65438 59950 65490
rect 60002 65438 60004 65490
rect 59948 65426 60004 65438
rect 60508 66164 60564 66174
rect 60508 64820 60564 66108
rect 60620 66050 60676 66062
rect 60620 65998 60622 66050
rect 60674 65998 60676 66050
rect 60620 65604 60676 65998
rect 60732 65604 60788 65614
rect 60620 65602 60788 65604
rect 60620 65550 60734 65602
rect 60786 65550 60788 65602
rect 60620 65548 60788 65550
rect 60732 65538 60788 65548
rect 60844 65044 60900 70588
rect 60956 70084 61012 71148
rect 61516 70978 61572 70990
rect 61516 70926 61518 70978
rect 61570 70926 61572 70978
rect 61516 70420 61572 70926
rect 61516 70354 61572 70364
rect 60956 70018 61012 70028
rect 61292 70082 61348 70094
rect 61292 70030 61294 70082
rect 61346 70030 61348 70082
rect 61180 68852 61236 68862
rect 61292 68852 61348 70030
rect 61180 68850 61348 68852
rect 61180 68798 61182 68850
rect 61234 68798 61348 68850
rect 61180 68796 61348 68798
rect 61180 68786 61236 68796
rect 61516 68628 61572 68638
rect 61516 68534 61572 68572
rect 61516 67732 61572 67742
rect 61516 67638 61572 67676
rect 61628 67508 61684 77644
rect 62076 77252 62132 77262
rect 62076 77158 62132 77196
rect 62636 75796 62692 78542
rect 62972 78596 63028 78606
rect 62972 77924 63028 78540
rect 63420 78372 63476 78382
rect 63420 78258 63476 78316
rect 63420 78206 63422 78258
rect 63474 78206 63476 78258
rect 63420 78194 63476 78206
rect 62972 77922 63140 77924
rect 62972 77870 62974 77922
rect 63026 77870 63140 77922
rect 62972 77868 63140 77870
rect 62972 77858 63028 77868
rect 63084 77364 63140 77868
rect 63084 77298 63140 77308
rect 62300 75740 62692 75796
rect 62972 77252 63028 77262
rect 62972 75796 63028 77196
rect 63532 76692 63588 76702
rect 63532 76598 63588 76636
rect 63868 76356 63924 76366
rect 63868 76262 63924 76300
rect 63980 76020 64036 78764
rect 64316 78754 64372 78764
rect 64316 77140 64372 77150
rect 64428 77140 64484 80108
rect 64764 80098 64820 80108
rect 65660 79604 65716 84476
rect 65772 84438 65828 84476
rect 65884 84308 65940 85036
rect 66220 84868 66276 84878
rect 66220 84774 66276 84812
rect 66332 84308 66388 84318
rect 65884 84306 66388 84308
rect 65884 84254 66334 84306
rect 66386 84254 66388 84306
rect 65884 84252 66388 84254
rect 65916 83916 66180 83926
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 65916 83850 66180 83860
rect 65916 82348 66180 82358
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 65916 82282 66180 82292
rect 65772 81396 65828 81406
rect 65772 80386 65828 81340
rect 66332 81396 66388 84252
rect 66444 84308 66500 85820
rect 67228 85876 67284 85886
rect 66556 85090 66612 85102
rect 66556 85038 66558 85090
rect 66610 85038 66612 85090
rect 66556 84532 66612 85038
rect 67116 85090 67172 85102
rect 67116 85038 67118 85090
rect 67170 85038 67172 85090
rect 67116 84980 67172 85038
rect 67116 84914 67172 84924
rect 67228 84978 67284 85820
rect 67452 85764 67508 87276
rect 68124 87330 68180 87342
rect 68124 87278 68126 87330
rect 68178 87278 68180 87330
rect 68124 86548 68180 87278
rect 68236 87332 68292 88958
rect 68908 88900 68964 88910
rect 70476 88900 70532 88910
rect 68908 88898 69412 88900
rect 68908 88846 68910 88898
rect 68962 88846 69412 88898
rect 68908 88844 69412 88846
rect 68908 88834 68964 88844
rect 68236 87266 68292 87276
rect 69244 86660 69300 86670
rect 68236 86548 68292 86558
rect 68124 86546 68292 86548
rect 68124 86494 68238 86546
rect 68290 86494 68292 86546
rect 68124 86492 68292 86494
rect 68236 86482 68292 86492
rect 68572 86548 68628 86558
rect 68572 86454 68628 86492
rect 67452 85698 67508 85708
rect 68348 86436 68404 86446
rect 68348 85090 68404 86380
rect 68348 85038 68350 85090
rect 68402 85038 68404 85090
rect 68348 85026 68404 85038
rect 67228 84926 67230 84978
rect 67282 84926 67284 84978
rect 67228 84914 67284 84926
rect 67340 84980 67396 84990
rect 66556 84466 66612 84476
rect 67116 84420 67172 84430
rect 67116 84326 67172 84364
rect 66444 84242 66500 84252
rect 67340 84084 67396 84924
rect 68012 84866 68068 84878
rect 68012 84814 68014 84866
rect 68066 84814 68068 84866
rect 68012 84420 68068 84814
rect 68012 84354 68068 84364
rect 69244 84194 69300 86604
rect 69244 84142 69246 84194
rect 69298 84142 69300 84194
rect 67340 84018 67396 84028
rect 67676 84084 67732 84094
rect 67676 83634 67732 84028
rect 67676 83582 67678 83634
rect 67730 83582 67732 83634
rect 67676 83570 67732 83582
rect 68684 82292 68740 82302
rect 66332 81330 66388 81340
rect 68012 81842 68068 81854
rect 68012 81790 68014 81842
rect 68066 81790 68068 81842
rect 66332 81058 66388 81070
rect 66332 81006 66334 81058
rect 66386 81006 66388 81058
rect 65916 80780 66180 80790
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 65916 80714 66180 80724
rect 65772 80334 65774 80386
rect 65826 80334 65828 80386
rect 65772 80322 65828 80334
rect 66332 79716 66388 81006
rect 68012 80388 68068 81790
rect 68124 81732 68180 81742
rect 68124 81730 68292 81732
rect 68124 81678 68126 81730
rect 68178 81678 68292 81730
rect 68124 81676 68292 81678
rect 68124 81666 68180 81676
rect 68012 80322 68068 80332
rect 68124 81060 68180 81070
rect 66444 80276 66500 80286
rect 66444 80274 66612 80276
rect 66444 80222 66446 80274
rect 66498 80222 66612 80274
rect 66444 80220 66612 80222
rect 66444 80210 66500 80220
rect 66444 79716 66500 79726
rect 66332 79660 66444 79716
rect 66444 79584 66500 79660
rect 65660 79538 65716 79548
rect 65916 79212 66180 79222
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 65916 79146 66180 79156
rect 66332 78932 66388 78942
rect 65100 78708 65156 78718
rect 65100 78706 65380 78708
rect 65100 78654 65102 78706
rect 65154 78654 65380 78706
rect 65100 78652 65380 78654
rect 65100 78642 65156 78652
rect 65324 78258 65380 78652
rect 65324 78206 65326 78258
rect 65378 78206 65380 78258
rect 65324 78194 65380 78206
rect 66332 78258 66388 78876
rect 66556 78820 66612 80220
rect 67452 79714 67508 79726
rect 67452 79662 67454 79714
rect 67506 79662 67508 79714
rect 66780 79602 66836 79614
rect 66780 79550 66782 79602
rect 66834 79550 66836 79602
rect 66780 79492 66836 79550
rect 66780 79426 66836 79436
rect 67228 79602 67284 79614
rect 67228 79550 67230 79602
rect 67282 79550 67284 79602
rect 67228 78932 67284 79550
rect 67228 78800 67284 78876
rect 66556 78754 66612 78764
rect 66332 78206 66334 78258
rect 66386 78206 66388 78258
rect 66332 78194 66388 78206
rect 64316 77138 64484 77140
rect 64316 77086 64318 77138
rect 64370 77086 64484 77138
rect 64316 77084 64484 77086
rect 65548 78146 65604 78158
rect 65548 78094 65550 78146
rect 65602 78094 65604 78146
rect 62188 75458 62244 75470
rect 62188 75406 62190 75458
rect 62242 75406 62244 75458
rect 61852 74114 61908 74126
rect 61852 74062 61854 74114
rect 61906 74062 61908 74114
rect 61852 74004 61908 74062
rect 61852 73938 61908 73948
rect 62188 73442 62244 75406
rect 62188 73390 62190 73442
rect 62242 73390 62244 73442
rect 62188 73378 62244 73390
rect 62076 73220 62132 73230
rect 62076 72770 62132 73164
rect 62076 72718 62078 72770
rect 62130 72718 62132 72770
rect 62076 72706 62132 72718
rect 62300 72660 62356 75740
rect 62972 75664 63028 75740
rect 63756 75964 64148 76020
rect 63756 75682 63812 75964
rect 63756 75630 63758 75682
rect 63810 75630 63812 75682
rect 63756 75618 63812 75630
rect 63868 75796 63924 75806
rect 62524 75570 62580 75582
rect 62524 75518 62526 75570
rect 62578 75518 62580 75570
rect 62412 74114 62468 74126
rect 62412 74062 62414 74114
rect 62466 74062 62468 74114
rect 62412 72772 62468 74062
rect 62524 72996 62580 75518
rect 63420 74786 63476 74798
rect 63420 74734 63422 74786
rect 63474 74734 63476 74786
rect 62636 74004 62692 74014
rect 63420 74004 63476 74734
rect 63868 74114 63924 75740
rect 63868 74062 63870 74114
rect 63922 74062 63924 74114
rect 63868 74050 63924 74062
rect 63980 74786 64036 74798
rect 63980 74734 63982 74786
rect 64034 74734 64036 74786
rect 62636 74002 63476 74004
rect 62636 73950 62638 74002
rect 62690 73950 63476 74002
rect 62636 73948 63476 73950
rect 62636 73938 62692 73948
rect 63420 73892 63700 73948
rect 62524 72930 62580 72940
rect 62412 72716 62692 72772
rect 62300 72604 62468 72660
rect 61740 72548 61796 72558
rect 61740 72454 61796 72492
rect 62188 71092 62244 71102
rect 62188 70998 62244 71036
rect 62188 68628 62244 68638
rect 62188 68534 62244 68572
rect 62300 68516 62356 68526
rect 61852 68404 61908 68414
rect 61852 68066 61908 68348
rect 61852 68014 61854 68066
rect 61906 68014 61908 68066
rect 61852 68002 61908 68014
rect 60844 64978 60900 64988
rect 61292 67452 61684 67508
rect 62300 67842 62356 68460
rect 62412 68404 62468 72604
rect 62636 72548 62692 72716
rect 62748 72548 62804 72558
rect 62636 72546 62804 72548
rect 62636 72494 62750 72546
rect 62802 72494 62804 72546
rect 62636 72492 62804 72494
rect 62748 72212 62804 72492
rect 62748 72146 62804 72156
rect 62860 72434 62916 72446
rect 62860 72382 62862 72434
rect 62914 72382 62916 72434
rect 62748 71762 62804 71774
rect 62748 71710 62750 71762
rect 62802 71710 62804 71762
rect 62748 71652 62804 71710
rect 62748 71586 62804 71596
rect 62860 71092 62916 72382
rect 63644 72434 63700 73892
rect 63644 72382 63646 72434
rect 63698 72382 63700 72434
rect 63644 72370 63700 72382
rect 63644 72212 63700 72222
rect 63644 71986 63700 72156
rect 63980 72212 64036 74734
rect 64092 73556 64148 75964
rect 64316 74900 64372 77084
rect 65436 77028 65492 77038
rect 65548 77028 65604 78094
rect 65660 78036 65716 78046
rect 66108 78036 66164 78046
rect 65660 78034 66164 78036
rect 65660 77982 65662 78034
rect 65714 77982 66110 78034
rect 66162 77982 66164 78034
rect 65660 77980 66164 77982
rect 65660 77970 65716 77980
rect 66108 77970 66164 77980
rect 66444 78036 66500 78046
rect 66892 78036 66948 78046
rect 66444 78034 66948 78036
rect 66444 77982 66446 78034
rect 66498 77982 66894 78034
rect 66946 77982 66948 78034
rect 66444 77980 66948 77982
rect 66444 77970 66500 77980
rect 65916 77644 66180 77654
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 65916 77578 66180 77588
rect 66668 77028 66724 77980
rect 66892 77970 66948 77980
rect 65548 76972 66612 77028
rect 64540 76692 64596 76702
rect 64540 76598 64596 76636
rect 65436 76690 65492 76972
rect 65436 76638 65438 76690
rect 65490 76638 65492 76690
rect 65436 76626 65492 76638
rect 66556 76804 66612 76972
rect 66668 76962 66724 76972
rect 66556 76748 67060 76804
rect 64764 76580 64820 76590
rect 64764 76486 64820 76524
rect 66444 76580 66500 76590
rect 66444 76486 66500 76524
rect 66556 76578 66612 76748
rect 67004 76690 67060 76748
rect 67004 76638 67006 76690
rect 67058 76638 67060 76690
rect 67004 76626 67060 76638
rect 66556 76526 66558 76578
rect 66610 76526 66612 76578
rect 66556 76514 66612 76526
rect 66668 76580 66724 76590
rect 64316 74806 64372 74844
rect 64428 76466 64484 76478
rect 64428 76414 64430 76466
rect 64482 76414 64484 76466
rect 64428 76356 64484 76414
rect 64428 75124 64484 76300
rect 65772 76466 65828 76478
rect 65772 76414 65774 76466
rect 65826 76414 65828 76466
rect 64540 75796 64596 75806
rect 64540 75702 64596 75740
rect 64428 74228 64484 75068
rect 65436 75124 65492 75134
rect 65436 75030 65492 75068
rect 65772 75124 65828 76414
rect 66444 76242 66500 76254
rect 66444 76190 66446 76242
rect 66498 76190 66500 76242
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 66444 75796 66500 76190
rect 66444 75730 66500 75740
rect 66668 75794 66724 76524
rect 67228 76580 67284 76590
rect 67228 76486 67284 76524
rect 66668 75742 66670 75794
rect 66722 75742 66724 75794
rect 66668 75730 66724 75742
rect 66780 76468 66836 76478
rect 66220 75684 66276 75694
rect 66220 75124 66276 75628
rect 65772 75122 66276 75124
rect 65772 75070 66222 75122
rect 66274 75070 66276 75122
rect 65772 75068 66276 75070
rect 65772 75010 65828 75068
rect 66220 75058 66276 75068
rect 65772 74958 65774 75010
rect 65826 74958 65828 75010
rect 65772 74946 65828 74958
rect 66780 74900 66836 76412
rect 67340 76466 67396 76478
rect 67340 76414 67342 76466
rect 67394 76414 67396 76466
rect 66892 76244 66948 76254
rect 66892 75684 66948 76188
rect 67228 76020 67284 76030
rect 67116 75684 67172 75694
rect 66948 75682 67172 75684
rect 66948 75630 67118 75682
rect 67170 75630 67172 75682
rect 66948 75628 67172 75630
rect 66892 75552 66948 75628
rect 67116 75618 67172 75628
rect 67004 74900 67060 74910
rect 66780 74898 67060 74900
rect 66780 74846 67006 74898
rect 67058 74846 67060 74898
rect 66780 74844 67060 74846
rect 67004 74834 67060 74844
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 64428 74162 64484 74172
rect 64092 73490 64148 73500
rect 65324 73556 65380 73566
rect 65324 73462 65380 73500
rect 65548 73556 65604 73566
rect 64316 73220 64372 73230
rect 64316 73218 64484 73220
rect 64316 73166 64318 73218
rect 64370 73166 64484 73218
rect 64316 73164 64484 73166
rect 64316 73154 64372 73164
rect 64428 72546 64484 73164
rect 64764 72996 64820 73006
rect 64764 72770 64820 72940
rect 64764 72718 64766 72770
rect 64818 72718 64820 72770
rect 64764 72706 64820 72718
rect 64428 72494 64430 72546
rect 64482 72494 64484 72546
rect 63980 72146 64036 72156
rect 64204 72434 64260 72446
rect 64204 72382 64206 72434
rect 64258 72382 64260 72434
rect 64204 72212 64260 72382
rect 64428 72324 64484 72494
rect 64428 72258 64484 72268
rect 65324 72322 65380 72334
rect 65324 72270 65326 72322
rect 65378 72270 65380 72322
rect 64204 72146 64260 72156
rect 65324 72212 65380 72270
rect 63644 71934 63646 71986
rect 63698 71934 63700 71986
rect 63644 71922 63700 71934
rect 63196 71652 63252 71662
rect 63196 71558 63252 71596
rect 63756 71652 63812 71662
rect 62860 71026 62916 71036
rect 63308 71092 63364 71102
rect 62972 70420 63028 70430
rect 62412 68338 62468 68348
rect 62524 68402 62580 68414
rect 62524 68350 62526 68402
rect 62578 68350 62580 68402
rect 62524 68068 62580 68350
rect 62524 68002 62580 68012
rect 62300 67790 62302 67842
rect 62354 67790 62356 67842
rect 61292 64820 61348 67452
rect 61628 66276 61684 66286
rect 61964 66276 62020 66286
rect 61628 66182 61684 66220
rect 61852 66274 62020 66276
rect 61852 66222 61966 66274
rect 62018 66222 62020 66274
rect 61852 66220 62020 66222
rect 61852 65604 61908 66220
rect 61964 66210 62020 66220
rect 62300 66162 62356 67790
rect 62300 66110 62302 66162
rect 62354 66110 62356 66162
rect 62300 66098 62356 66110
rect 62636 67730 62692 67742
rect 62636 67678 62638 67730
rect 62690 67678 62692 67730
rect 62636 66946 62692 67678
rect 62972 67172 63028 70364
rect 63308 68738 63364 71036
rect 63308 68686 63310 68738
rect 63362 68686 63364 68738
rect 63308 68674 63364 68686
rect 63420 70082 63476 70094
rect 63420 70030 63422 70082
rect 63474 70030 63476 70082
rect 63196 68628 63252 68666
rect 63196 68562 63252 68572
rect 63196 68404 63252 68414
rect 63196 67954 63252 68348
rect 63420 68068 63476 70030
rect 63644 68852 63700 68862
rect 63420 68002 63476 68012
rect 63532 68628 63588 68638
rect 63196 67902 63198 67954
rect 63250 67902 63252 67954
rect 63196 67890 63252 67902
rect 63532 67284 63588 68572
rect 63308 67282 63588 67284
rect 63308 67230 63534 67282
rect 63586 67230 63588 67282
rect 63308 67228 63588 67230
rect 63084 67172 63140 67182
rect 62972 67170 63252 67172
rect 62972 67118 63086 67170
rect 63138 67118 63252 67170
rect 62972 67116 63252 67118
rect 63084 67106 63140 67116
rect 62636 66894 62638 66946
rect 62690 66894 62692 66946
rect 62636 66162 62692 66894
rect 62636 66110 62638 66162
rect 62690 66110 62692 66162
rect 62636 66098 62692 66110
rect 63196 65716 63252 67116
rect 63308 66386 63364 67228
rect 63532 67218 63588 67228
rect 63308 66334 63310 66386
rect 63362 66334 63364 66386
rect 63308 66322 63364 66334
rect 63308 65716 63364 65726
rect 63196 65714 63364 65716
rect 63196 65662 63310 65714
rect 63362 65662 63364 65714
rect 63196 65660 63364 65662
rect 63308 65650 63364 65660
rect 59836 64708 59892 64718
rect 59836 64614 59892 64652
rect 60508 64594 60564 64764
rect 60620 64818 61348 64820
rect 60620 64766 61294 64818
rect 61346 64766 61348 64818
rect 60620 64764 61348 64766
rect 60620 64706 60676 64764
rect 61292 64754 61348 64764
rect 61740 64820 61796 64830
rect 60620 64654 60622 64706
rect 60674 64654 60676 64706
rect 60620 64642 60676 64654
rect 60508 64542 60510 64594
rect 60562 64542 60564 64594
rect 60508 64530 60564 64542
rect 60284 64484 60340 64494
rect 60284 64390 60340 64428
rect 61740 64484 61796 64764
rect 61740 64418 61796 64428
rect 61628 64372 61684 64382
rect 61628 64146 61684 64316
rect 61852 64260 61908 65548
rect 62860 65604 62916 65614
rect 62860 65378 62916 65548
rect 62860 65326 62862 65378
rect 62914 65326 62916 65378
rect 62860 65314 62916 65326
rect 61628 64094 61630 64146
rect 61682 64094 61684 64146
rect 61628 64082 61684 64094
rect 61740 64204 61908 64260
rect 61964 64260 62020 64270
rect 59724 63870 59726 63922
rect 59778 63870 59780 63922
rect 59724 63858 59780 63870
rect 60508 63922 60564 63934
rect 60508 63870 60510 63922
rect 60562 63870 60564 63922
rect 59612 63086 59614 63138
rect 59666 63086 59668 63138
rect 59612 63074 59668 63086
rect 60396 63812 60452 63822
rect 60060 63026 60116 63038
rect 60060 62974 60062 63026
rect 60114 62974 60116 63026
rect 59836 62914 59892 62926
rect 59836 62862 59838 62914
rect 59890 62862 59892 62914
rect 59276 62804 59332 62814
rect 59276 62578 59332 62748
rect 59276 62526 59278 62578
rect 59330 62526 59332 62578
rect 59276 62514 59332 62526
rect 59500 62580 59556 62590
rect 59836 62580 59892 62862
rect 59500 62578 59892 62580
rect 59500 62526 59502 62578
rect 59554 62526 59892 62578
rect 59500 62524 59892 62526
rect 60060 62580 60116 62974
rect 59500 62514 59556 62524
rect 60060 62514 60116 62524
rect 60284 62804 60340 62814
rect 60284 62578 60340 62748
rect 60284 62526 60286 62578
rect 60338 62526 60340 62578
rect 60284 62514 60340 62526
rect 59164 62354 59220 62366
rect 59164 62302 59166 62354
rect 59218 62302 59220 62354
rect 59164 62188 59220 62302
rect 59948 62242 60004 62254
rect 59948 62190 59950 62242
rect 60002 62190 60004 62242
rect 59948 62188 60004 62190
rect 59164 62132 60340 62188
rect 58940 61518 58942 61570
rect 58994 61518 58996 61570
rect 58940 61506 58996 61518
rect 59164 61460 59220 61470
rect 59164 61366 59220 61404
rect 59276 61458 59332 61470
rect 59276 61406 59278 61458
rect 59330 61406 59332 61458
rect 59276 61348 59332 61406
rect 60172 61460 60228 61470
rect 60172 61366 60228 61404
rect 59276 61282 59332 61292
rect 59724 61348 59780 61358
rect 59724 61254 59780 61292
rect 58604 61068 58772 61124
rect 59724 61124 59780 61134
rect 60284 61124 60340 62132
rect 57372 60788 57428 60798
rect 57372 60676 57428 60732
rect 57820 60676 57876 60686
rect 57372 60674 57876 60676
rect 57372 60622 57374 60674
rect 57426 60622 57822 60674
rect 57874 60622 57876 60674
rect 57372 60620 57876 60622
rect 57260 60228 57316 60238
rect 57260 60134 57316 60172
rect 57260 59892 57316 59902
rect 57260 59798 57316 59836
rect 57372 59890 57428 60620
rect 57820 60610 57876 60620
rect 57372 59838 57374 59890
rect 57426 59838 57428 59890
rect 57372 59780 57428 59838
rect 57372 59714 57428 59724
rect 58044 59892 58100 59902
rect 57596 59332 57652 59342
rect 57596 59238 57652 59276
rect 57708 59220 57764 59230
rect 57708 59126 57764 59164
rect 57596 58994 57652 59006
rect 57596 58942 57598 58994
rect 57650 58942 57652 58994
rect 57260 58884 57316 58894
rect 57260 57764 57316 58828
rect 57596 58660 57652 58942
rect 57596 58212 57652 58604
rect 57932 58996 57988 59006
rect 57932 58324 57988 58940
rect 58044 58546 58100 59836
rect 58380 59892 58436 59902
rect 58380 59798 58436 59836
rect 58492 59890 58548 59902
rect 58492 59838 58494 59890
rect 58546 59838 58548 59890
rect 58156 59778 58212 59790
rect 58156 59726 58158 59778
rect 58210 59726 58212 59778
rect 58156 59668 58212 59726
rect 58492 59780 58548 59838
rect 58492 59714 58548 59724
rect 58156 59602 58212 59612
rect 58492 59556 58548 59566
rect 58156 59444 58212 59454
rect 58156 59350 58212 59388
rect 58044 58494 58046 58546
rect 58098 58494 58100 58546
rect 58044 58482 58100 58494
rect 58380 59330 58436 59342
rect 58380 59278 58382 59330
rect 58434 59278 58436 59330
rect 57932 58268 58100 58324
rect 57596 58156 57876 58212
rect 57260 57698 57316 57708
rect 57372 57876 57428 57886
rect 57372 57652 57428 57820
rect 57596 57764 57652 57774
rect 57372 57090 57428 57596
rect 57372 57038 57374 57090
rect 57426 57038 57428 57090
rect 57372 57026 57428 57038
rect 57484 57762 57652 57764
rect 57484 57710 57598 57762
rect 57650 57710 57652 57762
rect 57484 57708 57652 57710
rect 57484 57092 57540 57708
rect 57596 57698 57652 57708
rect 57708 57764 57764 57774
rect 57708 57670 57764 57708
rect 57484 57026 57540 57036
rect 57596 57426 57652 57438
rect 57596 57374 57598 57426
rect 57650 57374 57652 57426
rect 57484 56868 57540 56878
rect 57484 56774 57540 56812
rect 57372 56756 57428 56766
rect 57372 56662 57428 56700
rect 57596 56420 57652 57374
rect 57596 56354 57652 56364
rect 57372 56308 57428 56318
rect 57372 56214 57428 56252
rect 57596 56196 57652 56206
rect 57036 55234 57092 55244
rect 57484 56194 57652 56196
rect 57484 56142 57598 56194
rect 57650 56142 57652 56194
rect 57484 56140 57652 56142
rect 56700 54686 56702 54738
rect 56754 54686 56756 54738
rect 56700 54674 56756 54686
rect 57036 55074 57092 55086
rect 57036 55022 57038 55074
rect 57090 55022 57092 55074
rect 55692 54626 55748 54638
rect 55692 54574 55694 54626
rect 55746 54574 55748 54626
rect 55692 54516 55748 54574
rect 56476 54626 56532 54638
rect 56476 54574 56478 54626
rect 56530 54574 56532 54626
rect 55692 54450 55748 54460
rect 55804 54516 55860 54526
rect 56364 54516 56420 54526
rect 55804 54514 56420 54516
rect 55804 54462 55806 54514
rect 55858 54462 56366 54514
rect 56418 54462 56420 54514
rect 55804 54460 56420 54462
rect 55804 54450 55860 54460
rect 55580 51998 55582 52050
rect 55634 51998 55636 52050
rect 55580 51986 55636 51998
rect 56028 54292 56084 54302
rect 55356 51650 55412 51660
rect 55244 51436 55412 51492
rect 55244 51266 55300 51278
rect 55244 51214 55246 51266
rect 55298 51214 55300 51266
rect 55244 51154 55300 51214
rect 55244 51102 55246 51154
rect 55298 51102 55300 51154
rect 55244 51090 55300 51102
rect 55244 50596 55300 50606
rect 55132 50594 55300 50596
rect 55132 50542 55246 50594
rect 55298 50542 55300 50594
rect 55132 50540 55300 50542
rect 55244 50530 55300 50540
rect 54908 50428 55188 50484
rect 55132 50372 55188 50428
rect 55132 50316 55300 50372
rect 54460 48862 54462 48914
rect 54514 48862 54516 48914
rect 53900 48468 53956 48478
rect 53900 48374 53956 48412
rect 54124 48356 54180 48366
rect 54124 48262 54180 48300
rect 53564 48132 53620 48142
rect 53340 47124 53396 47134
rect 53340 46898 53396 47068
rect 53340 46846 53342 46898
rect 53394 46846 53396 46898
rect 53340 46834 53396 46846
rect 53564 46898 53620 48076
rect 53676 47124 53732 48188
rect 53676 47058 53732 47068
rect 54236 48242 54292 48254
rect 54236 48190 54238 48242
rect 54290 48190 54292 48242
rect 53564 46846 53566 46898
rect 53618 46846 53620 46898
rect 53564 46834 53620 46846
rect 53676 46900 53732 46910
rect 53676 46786 53732 46844
rect 54236 46900 54292 48190
rect 54236 46806 54292 46844
rect 53676 46734 53678 46786
rect 53730 46734 53732 46786
rect 53676 46722 53732 46734
rect 53228 46620 53620 46676
rect 52892 44994 53060 44996
rect 52892 44942 52894 44994
rect 52946 44942 53060 44994
rect 52892 44940 53060 44942
rect 53452 44994 53508 45006
rect 53452 44942 53454 44994
rect 53506 44942 53508 44994
rect 52332 44100 52388 44110
rect 52332 44006 52388 44044
rect 52892 43708 52948 44940
rect 52220 43650 52276 43662
rect 52220 43598 52222 43650
rect 52274 43598 52276 43650
rect 52220 43540 52276 43598
rect 52780 43652 52948 43708
rect 53228 44100 53284 44110
rect 53228 43708 53284 44044
rect 53452 43708 53508 44942
rect 53228 43652 53508 43708
rect 52780 43558 52836 43596
rect 52220 43474 52276 43484
rect 52332 43316 52388 43326
rect 52332 41076 52388 43260
rect 52668 42866 52724 42878
rect 52668 42814 52670 42866
rect 52722 42814 52724 42866
rect 52668 42084 52724 42814
rect 52668 42018 52724 42028
rect 52444 41860 52500 41870
rect 52444 41766 52500 41804
rect 53116 41746 53172 41758
rect 53116 41694 53118 41746
rect 53170 41694 53172 41746
rect 52556 41300 52612 41310
rect 52556 41186 52612 41244
rect 52556 41134 52558 41186
rect 52610 41134 52612 41186
rect 52556 41122 52612 41134
rect 53116 41188 53172 41694
rect 53228 41410 53284 43652
rect 53452 43540 53508 43550
rect 53340 43426 53396 43438
rect 53340 43374 53342 43426
rect 53394 43374 53396 43426
rect 53340 43316 53396 43374
rect 53340 43250 53396 43260
rect 53452 42866 53508 43484
rect 53452 42814 53454 42866
rect 53506 42814 53508 42866
rect 53452 42802 53508 42814
rect 53452 41860 53508 41870
rect 53452 41766 53508 41804
rect 53228 41358 53230 41410
rect 53282 41358 53284 41410
rect 53228 41300 53284 41358
rect 53340 41300 53396 41310
rect 53228 41298 53396 41300
rect 53228 41246 53342 41298
rect 53394 41246 53396 41298
rect 53228 41244 53396 41246
rect 53116 41122 53172 41132
rect 52332 39508 52388 41020
rect 53340 40514 53396 41244
rect 53340 40462 53342 40514
rect 53394 40462 53396 40514
rect 53340 39620 53396 40462
rect 53452 39620 53508 39630
rect 53340 39618 53508 39620
rect 53340 39566 53454 39618
rect 53506 39566 53508 39618
rect 53340 39564 53508 39566
rect 52332 39442 52388 39452
rect 52220 38948 52276 38958
rect 53004 38948 53060 38958
rect 52108 38946 52276 38948
rect 52108 38894 52222 38946
rect 52274 38894 52276 38946
rect 52108 38892 52276 38894
rect 50652 38836 50708 38846
rect 51324 38836 51380 38846
rect 50652 38834 51380 38836
rect 50652 38782 50654 38834
rect 50706 38782 51326 38834
rect 51378 38782 51380 38834
rect 50652 38780 51380 38782
rect 50652 38770 50708 38780
rect 51324 38770 51380 38780
rect 51660 38612 51716 38622
rect 51436 38610 51716 38612
rect 51436 38558 51662 38610
rect 51714 38558 51716 38610
rect 51436 38556 51716 38558
rect 52220 38612 52276 38892
rect 52780 38946 53060 38948
rect 52780 38894 53006 38946
rect 53058 38894 53060 38946
rect 52780 38892 53060 38894
rect 52444 38836 52500 38846
rect 52780 38836 52836 38892
rect 53004 38882 53060 38892
rect 52444 38834 52836 38836
rect 52444 38782 52446 38834
rect 52498 38782 52836 38834
rect 52444 38780 52836 38782
rect 52444 38770 52500 38780
rect 52220 38556 52724 38612
rect 50540 38164 50596 38174
rect 50316 38162 50596 38164
rect 50316 38110 50542 38162
rect 50594 38110 50596 38162
rect 50316 38108 50596 38110
rect 50540 38098 50596 38108
rect 49756 38052 49812 38062
rect 49644 38050 49812 38052
rect 49644 37998 49758 38050
rect 49810 37998 49812 38050
rect 49644 37996 49812 37998
rect 49196 37826 49252 37838
rect 49196 37774 49198 37826
rect 49250 37774 49252 37826
rect 49196 37380 49252 37774
rect 49196 37314 49252 37324
rect 48972 36642 49028 36652
rect 49644 37266 49700 37996
rect 49756 37986 49812 37996
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50316 37380 50372 37390
rect 50316 37286 50372 37324
rect 49644 37214 49646 37266
rect 49698 37214 49700 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 49644 35700 49700 37214
rect 51436 37156 51492 38556
rect 51660 38546 51716 38556
rect 52668 38164 52724 38556
rect 52668 38032 52724 38108
rect 51100 36708 51156 36718
rect 51100 36614 51156 36652
rect 51436 36706 51492 37100
rect 52444 37156 52500 37166
rect 52444 37062 52500 37100
rect 51436 36654 51438 36706
rect 51490 36654 51492 36706
rect 51436 36642 51492 36654
rect 52220 36484 52276 36494
rect 52220 36390 52276 36428
rect 52780 36484 52836 38780
rect 53452 38836 53508 39564
rect 53452 38770 53508 38780
rect 52892 38724 52948 38734
rect 52892 37490 52948 38668
rect 53452 38164 53508 38174
rect 53452 38070 53508 38108
rect 52892 37438 52894 37490
rect 52946 37438 52948 37490
rect 52892 37426 52948 37438
rect 52780 36418 52836 36428
rect 53340 36484 53396 36494
rect 53340 36390 53396 36428
rect 52108 36372 52164 36382
rect 52108 36278 52164 36316
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 49980 35700 50036 35710
rect 49644 35698 50036 35700
rect 49644 35646 49982 35698
rect 50034 35646 50036 35698
rect 49644 35644 50036 35646
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 49868 34916 49924 34926
rect 49980 34916 50036 35644
rect 52892 35700 52948 35710
rect 53564 35700 53620 46620
rect 54460 46450 54516 48862
rect 54460 46398 54462 46450
rect 54514 46398 54516 46450
rect 54460 46386 54516 46398
rect 54684 49420 54852 49476
rect 55020 50260 55076 50270
rect 54124 45332 54180 45342
rect 53788 43540 53844 43550
rect 53788 43446 53844 43484
rect 54124 42754 54180 45276
rect 54348 43652 54404 43662
rect 54348 43558 54404 43596
rect 54124 42702 54126 42754
rect 54178 42702 54180 42754
rect 54124 42690 54180 42702
rect 54684 42196 54740 49420
rect 54908 48804 54964 48814
rect 54908 48710 54964 48748
rect 54796 48580 54852 48590
rect 54796 48020 54852 48524
rect 54908 48354 54964 48366
rect 54908 48302 54910 48354
rect 54962 48302 54964 48354
rect 54908 48244 54964 48302
rect 55020 48354 55076 50204
rect 55132 49924 55188 49934
rect 55132 48914 55188 49868
rect 55132 48862 55134 48914
rect 55186 48862 55188 48914
rect 55132 48850 55188 48862
rect 55244 48914 55300 50316
rect 55356 49812 55412 51436
rect 55692 51266 55748 51278
rect 55692 51214 55694 51266
rect 55746 51214 55748 51266
rect 55580 49924 55636 49934
rect 55580 49830 55636 49868
rect 55356 49810 55524 49812
rect 55356 49758 55358 49810
rect 55410 49758 55524 49810
rect 55356 49756 55524 49758
rect 55356 49680 55412 49756
rect 55244 48862 55246 48914
rect 55298 48862 55300 48914
rect 55020 48302 55022 48354
rect 55074 48302 55076 48354
rect 55020 48290 55076 48302
rect 54908 48178 54964 48188
rect 55244 48132 55300 48862
rect 55244 48066 55300 48076
rect 55468 48132 55524 49756
rect 55692 49028 55748 51214
rect 56028 51266 56084 54236
rect 56364 53732 56420 54460
rect 56476 54292 56532 54574
rect 56476 54226 56532 54236
rect 56364 53638 56420 53676
rect 56700 54068 56756 54078
rect 56700 53730 56756 54012
rect 56700 53678 56702 53730
rect 56754 53678 56756 53730
rect 56700 53666 56756 53678
rect 57036 53732 57092 55022
rect 57372 54402 57428 54414
rect 57372 54350 57374 54402
rect 57426 54350 57428 54402
rect 57372 54292 57428 54350
rect 57372 54226 57428 54236
rect 57484 54068 57540 56140
rect 57596 56130 57652 56140
rect 57708 56196 57764 56206
rect 57820 56196 57876 58156
rect 57932 57764 57988 57774
rect 57932 56866 57988 57708
rect 57932 56814 57934 56866
rect 57986 56814 57988 56866
rect 57932 56802 57988 56814
rect 57708 56194 57876 56196
rect 57708 56142 57710 56194
rect 57762 56142 57876 56194
rect 57708 56140 57876 56142
rect 57708 56130 57764 56140
rect 57484 54002 57540 54012
rect 57820 54402 57876 54414
rect 57820 54350 57822 54402
rect 57874 54350 57876 54402
rect 57036 53666 57092 53676
rect 57484 53732 57540 53742
rect 57484 53638 57540 53676
rect 57820 53732 57876 54350
rect 57820 53666 57876 53676
rect 56476 53508 56532 53518
rect 56476 53414 56532 53452
rect 57036 53508 57092 53518
rect 57148 53508 57204 53518
rect 57092 53506 57204 53508
rect 57092 53454 57150 53506
rect 57202 53454 57204 53506
rect 57092 53452 57204 53454
rect 56588 52276 56644 52286
rect 56252 52162 56308 52174
rect 56252 52110 56254 52162
rect 56306 52110 56308 52162
rect 56252 51492 56308 52110
rect 56588 52162 56644 52220
rect 56588 52110 56590 52162
rect 56642 52110 56644 52162
rect 56588 52098 56644 52110
rect 56252 51426 56308 51436
rect 56924 51492 56980 51502
rect 56028 51214 56030 51266
rect 56082 51214 56084 51266
rect 56028 49924 56084 51214
rect 56364 50820 56420 50830
rect 56364 50594 56420 50764
rect 56364 50542 56366 50594
rect 56418 50542 56420 50594
rect 56364 50530 56420 50542
rect 56812 50708 56868 50718
rect 56028 49858 56084 49868
rect 56476 50036 56532 50046
rect 56476 49810 56532 49980
rect 56700 50036 56756 50046
rect 56700 49942 56756 49980
rect 56476 49758 56478 49810
rect 56530 49758 56532 49810
rect 56476 49588 56532 49758
rect 56476 49522 56532 49532
rect 55804 49028 55860 49038
rect 55692 49026 55860 49028
rect 55692 48974 55806 49026
rect 55858 48974 55860 49026
rect 55692 48972 55860 48974
rect 55692 48132 55748 48142
rect 55468 48130 55636 48132
rect 55468 48078 55470 48130
rect 55522 48078 55636 48130
rect 55468 48076 55636 48078
rect 55468 48066 55524 48076
rect 54908 48020 54964 48030
rect 54796 48018 54964 48020
rect 54796 47966 54910 48018
rect 54962 47966 54964 48018
rect 54796 47964 54964 47966
rect 54908 47954 54964 47964
rect 55244 47796 55300 47806
rect 54908 47460 54964 47470
rect 54908 47366 54964 47404
rect 55244 46900 55300 47740
rect 55244 46768 55300 46844
rect 54796 46562 54852 46574
rect 54796 46510 54798 46562
rect 54850 46510 54852 46562
rect 54796 46450 54852 46510
rect 54796 46398 54798 46450
rect 54850 46398 54852 46450
rect 54796 46386 54852 46398
rect 55468 46450 55524 46462
rect 55468 46398 55470 46450
rect 55522 46398 55524 46450
rect 55468 45890 55524 46398
rect 55468 45838 55470 45890
rect 55522 45838 55524 45890
rect 55468 45332 55524 45838
rect 55356 45276 55468 45332
rect 55356 44322 55412 45276
rect 55468 45200 55524 45276
rect 55356 44270 55358 44322
rect 55410 44270 55412 44322
rect 55356 44258 55412 44270
rect 55580 43708 55636 48076
rect 55692 46898 55748 48076
rect 55804 47572 55860 48972
rect 56588 48914 56644 48926
rect 56588 48862 56590 48914
rect 56642 48862 56644 48914
rect 56588 48468 56644 48862
rect 56588 48402 56644 48412
rect 56476 48356 56532 48366
rect 56476 48262 56532 48300
rect 56252 48242 56308 48254
rect 56252 48190 56254 48242
rect 56306 48190 56308 48242
rect 55804 47570 56084 47572
rect 55804 47518 55806 47570
rect 55858 47518 56084 47570
rect 55804 47516 56084 47518
rect 55804 47506 55860 47516
rect 55692 46846 55694 46898
rect 55746 46846 55748 46898
rect 55692 46834 55748 46846
rect 56028 46898 56084 47516
rect 56028 46846 56030 46898
rect 56082 46846 56084 46898
rect 56028 46450 56084 46846
rect 56028 46398 56030 46450
rect 56082 46398 56084 46450
rect 56028 46386 56084 46398
rect 56140 46004 56196 46014
rect 56252 46004 56308 48190
rect 56588 48244 56644 48254
rect 56588 48150 56644 48188
rect 56140 46002 56308 46004
rect 56140 45950 56142 46002
rect 56194 45950 56308 46002
rect 56140 45948 56308 45950
rect 56140 45938 56196 45948
rect 56700 45332 56756 45342
rect 56252 45220 56308 45230
rect 56028 45218 56308 45220
rect 56028 45166 56254 45218
rect 56306 45166 56308 45218
rect 56028 45164 56308 45166
rect 56028 44434 56084 45164
rect 56252 45154 56308 45164
rect 56028 44382 56030 44434
rect 56082 44382 56084 44434
rect 56028 44370 56084 44382
rect 56588 45106 56644 45118
rect 56588 45054 56590 45106
rect 56642 45054 56644 45106
rect 55020 43652 55076 43662
rect 55580 43652 55748 43708
rect 54796 43650 55076 43652
rect 54796 43598 55022 43650
rect 55074 43598 55076 43650
rect 54796 43596 55076 43598
rect 54796 42866 54852 43596
rect 55020 43586 55076 43596
rect 54796 42814 54798 42866
rect 54850 42814 54852 42866
rect 54796 42802 54852 42814
rect 55356 43538 55412 43550
rect 55356 43486 55358 43538
rect 55410 43486 55412 43538
rect 54796 42196 54852 42206
rect 54684 42194 54852 42196
rect 54684 42142 54798 42194
rect 54850 42142 54852 42194
rect 54684 42140 54852 42142
rect 54124 42084 54180 42094
rect 54124 41990 54180 42028
rect 54684 42084 54740 42140
rect 54796 42130 54852 42140
rect 54684 42018 54740 42028
rect 54236 41970 54292 41982
rect 54236 41918 54238 41970
rect 54290 41918 54292 41970
rect 53788 41410 53844 41422
rect 53788 41358 53790 41410
rect 53842 41358 53844 41410
rect 53788 41298 53844 41358
rect 53788 41246 53790 41298
rect 53842 41246 53844 41298
rect 53788 41234 53844 41246
rect 54236 41300 54292 41918
rect 55356 41972 55412 43486
rect 55468 41972 55524 41982
rect 55356 41970 55524 41972
rect 55356 41918 55470 41970
rect 55522 41918 55524 41970
rect 55356 41916 55524 41918
rect 55468 41906 55524 41916
rect 54236 41206 54292 41244
rect 55132 41300 55188 41310
rect 55132 41206 55188 41244
rect 54684 41076 54740 41086
rect 54684 40982 54740 41020
rect 55580 40404 55636 40414
rect 55580 40310 55636 40348
rect 53676 39508 53732 39518
rect 53676 36596 53732 39452
rect 55468 39394 55524 39406
rect 55468 39342 55470 39394
rect 55522 39342 55524 39394
rect 54572 38948 54628 38958
rect 54572 38854 54628 38892
rect 55468 38948 55524 39342
rect 55468 38882 55524 38892
rect 53788 38836 53844 38846
rect 53788 38162 53844 38780
rect 53788 38110 53790 38162
rect 53842 38110 53844 38162
rect 53788 38098 53844 38110
rect 55692 38052 55748 43652
rect 56588 43652 56644 45054
rect 56588 43586 56644 43596
rect 56700 44436 56756 45276
rect 56700 43650 56756 44380
rect 56700 43598 56702 43650
rect 56754 43598 56756 43650
rect 56700 43586 56756 43598
rect 56812 42868 56868 50652
rect 56924 50594 56980 51436
rect 56924 50542 56926 50594
rect 56978 50542 56980 50594
rect 56924 50530 56980 50542
rect 57036 50036 57092 53452
rect 57148 53442 57204 53452
rect 57596 52164 57652 52174
rect 57596 52070 57652 52108
rect 57372 51604 57428 51614
rect 58044 51604 58100 58268
rect 58380 57876 58436 59278
rect 58492 59330 58548 59500
rect 58492 59278 58494 59330
rect 58546 59278 58548 59330
rect 58492 59266 58548 59278
rect 58492 58436 58548 58446
rect 58492 58342 58548 58380
rect 58380 57810 58436 57820
rect 58268 56756 58324 56766
rect 58268 56662 58324 56700
rect 58156 56644 58212 56654
rect 58156 56550 58212 56588
rect 58156 56084 58212 56094
rect 58156 55970 58212 56028
rect 58156 55918 58158 55970
rect 58210 55918 58212 55970
rect 58156 55524 58212 55918
rect 58604 55468 58660 61068
rect 58940 59778 58996 59790
rect 58940 59726 58942 59778
rect 58994 59726 58996 59778
rect 58940 59668 58996 59726
rect 58940 59602 58996 59612
rect 58940 59220 58996 59230
rect 58940 59106 58996 59164
rect 58940 59054 58942 59106
rect 58994 59054 58996 59106
rect 58716 56756 58772 56766
rect 58716 56644 58772 56700
rect 58940 56644 58996 59054
rect 59612 59218 59668 59230
rect 59612 59166 59614 59218
rect 59666 59166 59668 59218
rect 59612 58436 59668 59166
rect 59612 58370 59668 58380
rect 59164 56644 59220 56654
rect 58716 56642 59220 56644
rect 58716 56590 58718 56642
rect 58770 56590 59166 56642
rect 59218 56590 59220 56642
rect 58716 56588 59220 56590
rect 58716 56578 58772 56588
rect 59164 56084 59220 56588
rect 59164 56018 59220 56028
rect 59724 55468 59780 61068
rect 60172 61068 60340 61124
rect 60396 61124 60452 63756
rect 59836 58436 59892 58446
rect 59836 58342 59892 58380
rect 58156 55412 58212 55468
rect 58156 55346 58212 55356
rect 58492 55412 58660 55468
rect 59612 55412 59780 55468
rect 58268 51940 58324 51950
rect 58268 51846 58324 51884
rect 57372 51602 58100 51604
rect 57372 51550 57374 51602
rect 57426 51550 58100 51602
rect 57372 51548 58100 51550
rect 57372 51538 57428 51548
rect 58044 51378 58100 51548
rect 58044 51326 58046 51378
rect 58098 51326 58100 51378
rect 58044 51314 58100 51326
rect 57372 51156 57428 51166
rect 57372 50370 57428 51100
rect 58380 50708 58436 50718
rect 58380 50614 58436 50652
rect 57484 50596 57540 50606
rect 57484 50502 57540 50540
rect 58044 50596 58100 50606
rect 58044 50502 58100 50540
rect 57372 50318 57374 50370
rect 57426 50318 57428 50370
rect 57372 50306 57428 50318
rect 57596 50484 57652 50494
rect 57036 48804 57092 49980
rect 57596 50034 57652 50428
rect 57596 49982 57598 50034
rect 57650 49982 57652 50034
rect 57596 49970 57652 49982
rect 57484 49812 57540 49822
rect 57484 49718 57540 49756
rect 57820 49812 57876 49822
rect 57820 49810 58100 49812
rect 57820 49758 57822 49810
rect 57874 49758 58100 49810
rect 57820 49756 58100 49758
rect 57820 49746 57876 49756
rect 57036 48738 57092 48748
rect 57484 49588 57540 49598
rect 57372 48356 57428 48366
rect 57372 48262 57428 48300
rect 57484 48132 57540 49532
rect 57372 48076 57540 48132
rect 57596 48804 57652 48814
rect 57596 48466 57652 48748
rect 57596 48414 57598 48466
rect 57650 48414 57652 48466
rect 57372 43708 57428 48076
rect 57484 46900 57540 46910
rect 57596 46900 57652 48414
rect 58044 48356 58100 49756
rect 58156 49698 58212 49710
rect 58156 49646 58158 49698
rect 58210 49646 58212 49698
rect 58156 49588 58212 49646
rect 58156 49522 58212 49532
rect 58268 48356 58324 48366
rect 58044 48354 58324 48356
rect 58044 48302 58270 48354
rect 58322 48302 58324 48354
rect 58044 48300 58324 48302
rect 58268 48290 58324 48300
rect 58380 48354 58436 48366
rect 58380 48302 58382 48354
rect 58434 48302 58436 48354
rect 57708 48242 57764 48254
rect 57708 48190 57710 48242
rect 57762 48190 57764 48242
rect 57708 48132 57764 48190
rect 58380 48244 58436 48302
rect 58380 48178 58436 48188
rect 57708 48066 57764 48076
rect 57484 46898 57652 46900
rect 57484 46846 57486 46898
rect 57538 46846 57652 46898
rect 57484 46844 57652 46846
rect 58268 47124 58324 47134
rect 58492 47124 58548 55412
rect 59276 54402 59332 54414
rect 59276 54350 59278 54402
rect 59330 54350 59332 54402
rect 59276 54292 59332 54350
rect 59276 54226 59332 54236
rect 58716 52162 58772 52174
rect 58716 52110 58718 52162
rect 58770 52110 58772 52162
rect 58716 51604 58772 52110
rect 58716 51538 58772 51548
rect 58940 51940 58996 51950
rect 58716 51380 58772 51390
rect 58716 50484 58772 51324
rect 58604 49812 58660 49822
rect 58604 49698 58660 49756
rect 58604 49646 58606 49698
rect 58658 49646 58660 49698
rect 58604 49252 58660 49646
rect 58604 49186 58660 49196
rect 58716 49138 58772 50428
rect 58716 49086 58718 49138
rect 58770 49086 58772 49138
rect 58716 49074 58772 49086
rect 58828 50820 58884 50830
rect 58604 48468 58660 48478
rect 58604 48374 58660 48412
rect 57484 46834 57540 46844
rect 58268 46002 58324 47068
rect 58268 45950 58270 46002
rect 58322 45950 58324 46002
rect 58268 45938 58324 45950
rect 58380 47068 58548 47124
rect 58156 44548 58212 44558
rect 58156 44434 58212 44492
rect 58156 44382 58158 44434
rect 58210 44382 58212 44434
rect 58156 44370 58212 44382
rect 57372 43652 57540 43708
rect 56924 42868 56980 42878
rect 56588 42866 56980 42868
rect 56588 42814 56926 42866
rect 56978 42814 56980 42866
rect 56588 42812 56980 42814
rect 56588 42082 56644 42812
rect 56924 42802 56980 42812
rect 56588 42030 56590 42082
rect 56642 42030 56644 42082
rect 56476 41972 56532 41982
rect 56476 41878 56532 41916
rect 55804 41748 55860 41758
rect 55804 41746 56532 41748
rect 55804 41694 55806 41746
rect 55858 41694 56532 41746
rect 55804 41692 56532 41694
rect 55804 41682 55860 41692
rect 56028 40404 56084 40414
rect 56028 40310 56084 40348
rect 55804 39508 55860 39518
rect 56476 39508 56532 41692
rect 56588 41298 56644 42030
rect 57036 41972 57092 41982
rect 56588 41246 56590 41298
rect 56642 41246 56644 41298
rect 56588 41234 56644 41246
rect 56924 41860 56980 41870
rect 56924 41412 56980 41804
rect 56924 41298 56980 41356
rect 56924 41246 56926 41298
rect 56978 41246 56980 41298
rect 56924 41234 56980 41246
rect 57036 40404 57092 41916
rect 55804 39506 56420 39508
rect 55804 39454 55806 39506
rect 55858 39454 56420 39506
rect 55804 39452 56420 39454
rect 56476 39452 56756 39508
rect 55804 39442 55860 39452
rect 56364 38274 56420 39452
rect 56364 38222 56366 38274
rect 56418 38222 56420 38274
rect 56364 38210 56420 38222
rect 56700 38722 56756 39452
rect 56700 38670 56702 38722
rect 56754 38670 56756 38722
rect 56700 38274 56756 38670
rect 56700 38222 56702 38274
rect 56754 38222 56756 38274
rect 56700 38210 56756 38222
rect 55580 37996 55748 38052
rect 53788 36596 53844 36606
rect 53676 36594 53844 36596
rect 53676 36542 53790 36594
rect 53842 36542 53844 36594
rect 53676 36540 53844 36542
rect 53676 36372 53732 36540
rect 53788 36530 53844 36540
rect 54348 36596 54404 36606
rect 53676 36306 53732 36316
rect 54124 36484 54180 36494
rect 54124 35924 54180 36428
rect 54236 36260 54292 36270
rect 54348 36260 54404 36540
rect 55580 36596 55636 37996
rect 55580 36530 55636 36540
rect 55692 37828 55748 37838
rect 54236 36258 54404 36260
rect 54236 36206 54238 36258
rect 54290 36206 54404 36258
rect 54236 36204 54404 36206
rect 54236 36194 54292 36204
rect 54124 35810 54180 35868
rect 54124 35758 54126 35810
rect 54178 35758 54180 35810
rect 54124 35746 54180 35758
rect 50764 35588 50820 35598
rect 50764 35586 51044 35588
rect 50764 35534 50766 35586
rect 50818 35534 51044 35586
rect 50764 35532 51044 35534
rect 50764 35522 50820 35532
rect 49924 34860 50036 34916
rect 49868 34822 49924 34860
rect 50540 34804 50596 34814
rect 50540 34802 50932 34804
rect 50540 34750 50542 34802
rect 50594 34750 50932 34802
rect 50540 34748 50932 34750
rect 50540 34738 50596 34748
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50876 34020 50932 34748
rect 50988 34354 51044 35532
rect 52892 35586 52948 35644
rect 52892 35534 52894 35586
rect 52946 35534 52948 35586
rect 52892 35522 52948 35534
rect 53452 35644 53564 35700
rect 50988 34302 50990 34354
rect 51042 34302 51044 34354
rect 50988 34290 51044 34302
rect 51324 35476 51380 35486
rect 51324 34242 51380 35420
rect 52668 35364 52724 35374
rect 52668 35028 52724 35308
rect 51324 34190 51326 34242
rect 51378 34190 51380 34242
rect 51324 34178 51380 34190
rect 52332 35026 52724 35028
rect 52332 34974 52670 35026
rect 52722 34974 52724 35026
rect 52332 34972 52724 34974
rect 52332 34130 52388 34972
rect 52668 34962 52724 34972
rect 53452 35026 53508 35644
rect 53564 35634 53620 35644
rect 53564 35476 53620 35486
rect 53564 35382 53620 35420
rect 53900 35474 53956 35486
rect 53900 35422 53902 35474
rect 53954 35422 53956 35474
rect 53900 35364 53956 35422
rect 53900 35298 53956 35308
rect 53452 34974 53454 35026
rect 53506 34974 53508 35026
rect 53452 34962 53508 34974
rect 53676 34916 53732 34926
rect 53004 34804 53060 34814
rect 53004 34242 53060 34748
rect 53004 34190 53006 34242
rect 53058 34190 53060 34242
rect 53004 34178 53060 34190
rect 53676 34692 53732 34860
rect 54012 34804 54068 34814
rect 53788 34692 53844 34702
rect 53676 34690 53844 34692
rect 53676 34638 53790 34690
rect 53842 34638 53844 34690
rect 53676 34636 53844 34638
rect 52332 34078 52334 34130
rect 52386 34078 52388 34130
rect 52332 34066 52388 34078
rect 53116 34130 53172 34142
rect 53116 34078 53118 34130
rect 53170 34078 53172 34130
rect 50876 33964 51268 34020
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 51212 33236 51268 33964
rect 51996 33908 52052 33918
rect 51660 33906 52052 33908
rect 51660 33854 51998 33906
rect 52050 33854 52052 33906
rect 51660 33852 52052 33854
rect 51660 33346 51716 33852
rect 51996 33842 52052 33852
rect 53116 33460 53172 34078
rect 53116 33394 53172 33404
rect 53452 33460 53508 33470
rect 53676 33460 53732 34636
rect 53788 34626 53844 34636
rect 53900 34132 53956 34142
rect 53900 34038 53956 34076
rect 53452 33458 53732 33460
rect 53452 33406 53454 33458
rect 53506 33406 53732 33458
rect 53452 33404 53732 33406
rect 53788 33460 53844 33470
rect 53452 33394 53508 33404
rect 53788 33366 53844 33404
rect 51660 33294 51662 33346
rect 51714 33294 51716 33346
rect 51660 33282 51716 33294
rect 51324 33236 51380 33246
rect 51212 33234 51380 33236
rect 51212 33182 51326 33234
rect 51378 33182 51380 33234
rect 51212 33180 51380 33182
rect 51324 33170 51380 33180
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 53788 32788 53844 32798
rect 54012 32788 54068 34748
rect 53788 32786 54068 32788
rect 53788 32734 53790 32786
rect 53842 32734 54068 32786
rect 53788 32732 54068 32734
rect 54348 34802 54404 36204
rect 55244 35924 55300 35934
rect 55244 35830 55300 35868
rect 54460 35810 54516 35822
rect 54460 35758 54462 35810
rect 54514 35758 54516 35810
rect 54460 35700 54516 35758
rect 54460 35634 54516 35644
rect 54348 34750 54350 34802
rect 54402 34750 54404 34802
rect 53788 32722 53844 32732
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 18620 3444 18676 3454
rect 19068 3444 19124 3454
rect 18620 3442 19124 3444
rect 18620 3390 18622 3442
rect 18674 3390 19070 3442
rect 19122 3390 19124 3442
rect 18620 3388 19124 3390
rect 18620 3378 18676 3388
rect 14252 3266 14308 3276
rect 18844 800 18900 3388
rect 19068 3378 19124 3388
rect 31052 3444 31108 3454
rect 31500 3444 31556 3454
rect 31052 3442 31556 3444
rect 31052 3390 31054 3442
rect 31106 3390 31502 3442
rect 31554 3390 31556 3442
rect 31052 3388 31556 3390
rect 31052 3378 31108 3388
rect 19404 3332 19460 3342
rect 19404 3238 19460 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 31276 800 31332 3388
rect 31500 3378 31556 3388
rect 43708 3444 43764 3454
rect 31836 3330 31892 3342
rect 31836 3278 31838 3330
rect 31890 3278 31892 3330
rect 31836 2884 31892 3278
rect 31836 2818 31892 2828
rect 43708 800 43764 3388
rect 44268 3444 44324 3454
rect 44268 3350 44324 3388
rect 44940 3444 44996 3454
rect 44940 3350 44996 3388
rect 45276 3330 45332 3342
rect 45276 3278 45278 3330
rect 45330 3278 45332 3330
rect 45276 2772 45332 3278
rect 54348 3332 54404 34750
rect 54684 34804 54740 34814
rect 54684 34710 54740 34748
rect 55692 34804 55748 37772
rect 56700 37378 56756 37390
rect 56700 37326 56702 37378
rect 56754 37326 56756 37378
rect 56476 37268 56532 37278
rect 56476 37174 56532 37212
rect 56700 36596 56756 37326
rect 56812 36596 56868 36606
rect 56700 36594 56868 36596
rect 56700 36542 56814 36594
rect 56866 36542 56868 36594
rect 56700 36540 56868 36542
rect 56812 36530 56868 36540
rect 56140 36484 56196 36494
rect 56140 36482 56756 36484
rect 56140 36430 56142 36482
rect 56194 36430 56756 36482
rect 56140 36428 56756 36430
rect 56140 36418 56196 36428
rect 55692 34738 55748 34748
rect 56700 35922 56756 36428
rect 57036 36148 57092 40348
rect 57372 38050 57428 38062
rect 57372 37998 57374 38050
rect 57426 37998 57428 38050
rect 57260 37938 57316 37950
rect 57260 37886 57262 37938
rect 57314 37886 57316 37938
rect 57260 37828 57316 37886
rect 57260 37762 57316 37772
rect 57372 37716 57428 37998
rect 57372 37650 57428 37660
rect 56700 35870 56702 35922
rect 56754 35870 56756 35922
rect 56700 35028 56756 35870
rect 56700 34244 56756 34972
rect 56812 36092 57092 36148
rect 56812 34914 56868 36092
rect 57484 36036 57540 43652
rect 57596 43652 57652 43662
rect 57596 43558 57652 43596
rect 57932 43314 57988 43326
rect 57932 43262 57934 43314
rect 57986 43262 57988 43314
rect 57932 42868 57988 43262
rect 57932 42802 57988 42812
rect 57596 42754 57652 42766
rect 57596 42702 57598 42754
rect 57650 42702 57652 42754
rect 57596 41972 57652 42702
rect 58268 42644 58324 42654
rect 57596 41906 57652 41916
rect 57932 42642 58324 42644
rect 57932 42590 58270 42642
rect 58322 42590 58324 42642
rect 57932 42588 58324 42590
rect 57708 41188 57764 41198
rect 57708 41094 57764 41132
rect 57932 41074 57988 42588
rect 58268 42578 58324 42588
rect 57932 41022 57934 41074
rect 57986 41022 57988 41074
rect 57932 41010 57988 41022
rect 58156 40964 58212 40974
rect 58156 40402 58212 40908
rect 58156 40350 58158 40402
rect 58210 40350 58212 40402
rect 58044 37826 58100 37838
rect 58044 37774 58046 37826
rect 58098 37774 58100 37826
rect 58044 37716 58100 37774
rect 58156 37828 58212 40350
rect 58156 37762 58212 37772
rect 58044 37650 58100 37660
rect 57708 37268 57764 37278
rect 57708 37174 57764 37212
rect 58044 37044 58100 37054
rect 58044 37042 58212 37044
rect 58044 36990 58046 37042
rect 58098 36990 58212 37042
rect 58044 36988 58212 36990
rect 58044 36978 58100 36988
rect 57484 35980 57652 36036
rect 57484 35476 57540 35486
rect 57372 35028 57428 35038
rect 57372 34934 57428 34972
rect 56812 34862 56814 34914
rect 56866 34862 56868 34914
rect 56812 34850 56868 34862
rect 56700 34178 56756 34188
rect 54460 34132 54516 34142
rect 54460 33346 54516 34076
rect 54460 33294 54462 33346
rect 54514 33294 54516 33346
rect 54460 33282 54516 33294
rect 54572 34018 54628 34030
rect 54572 33966 54574 34018
rect 54626 33966 54628 34018
rect 54460 32788 54516 32798
rect 54572 32788 54628 33966
rect 56700 34020 56756 34030
rect 54460 32786 54628 32788
rect 54460 32734 54462 32786
rect 54514 32734 54628 32786
rect 54460 32732 54628 32734
rect 55244 33234 55300 33246
rect 55244 33182 55246 33234
rect 55298 33182 55300 33234
rect 54460 32722 54516 32732
rect 54796 32564 54852 32574
rect 54796 32470 54852 32508
rect 55244 31948 55300 33182
rect 56476 33236 56532 33246
rect 55916 33124 55972 33134
rect 55468 32564 55524 32574
rect 55468 32470 55524 32508
rect 55804 32564 55860 32574
rect 55804 32470 55860 32508
rect 55244 31892 55412 31948
rect 55356 31836 55636 31892
rect 55580 31666 55636 31836
rect 55916 31778 55972 33068
rect 56476 32562 56532 33180
rect 56588 32676 56644 32686
rect 56700 32676 56756 33964
rect 57484 34018 57540 35420
rect 57484 33966 57486 34018
rect 57538 33966 57540 34018
rect 57484 33954 57540 33966
rect 57372 33458 57428 33470
rect 57372 33406 57374 33458
rect 57426 33406 57428 33458
rect 57372 33348 57428 33406
rect 56588 32674 56756 32676
rect 56588 32622 56590 32674
rect 56642 32622 56756 32674
rect 56588 32620 56756 32622
rect 57036 33236 57092 33246
rect 56588 32610 56644 32620
rect 56476 32510 56478 32562
rect 56530 32510 56532 32562
rect 56476 32498 56532 32510
rect 57036 31890 57092 33180
rect 57372 32564 57428 33292
rect 57372 32498 57428 32508
rect 57596 32562 57652 35980
rect 58044 35812 58100 35822
rect 58044 35718 58100 35756
rect 58156 35476 58212 36988
rect 58156 35410 58212 35420
rect 58268 34132 58324 34142
rect 57932 34020 57988 34030
rect 57820 32788 57876 32798
rect 57820 32694 57876 32732
rect 57596 32510 57598 32562
rect 57650 32510 57652 32562
rect 57596 31948 57652 32510
rect 57036 31838 57038 31890
rect 57090 31838 57092 31890
rect 57036 31826 57092 31838
rect 57372 31892 57652 31948
rect 55916 31726 55918 31778
rect 55970 31726 55972 31778
rect 55916 31714 55972 31726
rect 55580 31614 55582 31666
rect 55634 31614 55636 31666
rect 55580 31602 55636 31614
rect 57372 31554 57428 31892
rect 57932 31890 57988 33964
rect 58044 33124 58100 33134
rect 58044 33030 58100 33068
rect 58268 32788 58324 34076
rect 58380 34020 58436 47068
rect 58716 45668 58772 45678
rect 58604 45666 58772 45668
rect 58604 45614 58718 45666
rect 58770 45614 58772 45666
rect 58604 45612 58772 45614
rect 58492 44548 58548 44558
rect 58492 43650 58548 44492
rect 58604 44436 58660 45612
rect 58716 45602 58772 45612
rect 58828 44548 58884 50764
rect 58940 50706 58996 51884
rect 59388 51492 59444 51502
rect 59164 51378 59220 51390
rect 59164 51326 59166 51378
rect 59218 51326 59220 51378
rect 59164 51044 59220 51326
rect 59164 50978 59220 50988
rect 58940 50654 58942 50706
rect 58994 50654 58996 50706
rect 58940 50596 58996 50654
rect 59388 50706 59444 51436
rect 59388 50654 59390 50706
rect 59442 50654 59444 50706
rect 59388 50642 59444 50654
rect 58940 50530 58996 50540
rect 59164 48356 59220 48366
rect 59052 48354 59220 48356
rect 59052 48302 59166 48354
rect 59218 48302 59220 48354
rect 59052 48300 59220 48302
rect 58940 48244 58996 48254
rect 58940 48150 58996 48188
rect 59052 47124 59108 48300
rect 59164 48290 59220 48300
rect 59276 48242 59332 48254
rect 59276 48190 59278 48242
rect 59330 48190 59332 48242
rect 59276 47796 59332 48190
rect 59276 47236 59332 47740
rect 59500 47236 59556 47246
rect 59276 47234 59556 47236
rect 59276 47182 59502 47234
rect 59554 47182 59556 47234
rect 59276 47180 59556 47182
rect 59052 47058 59108 47068
rect 59500 47124 59556 47180
rect 59500 47058 59556 47068
rect 58828 44482 58884 44492
rect 59276 44548 59332 44558
rect 58604 44342 58660 44380
rect 59276 44434 59332 44492
rect 59276 44382 59278 44434
rect 59330 44382 59332 44434
rect 59276 44370 59332 44382
rect 59612 43876 59668 55412
rect 59724 54740 59780 54750
rect 59724 54646 59780 54684
rect 59948 54626 60004 54638
rect 59948 54574 59950 54626
rect 60002 54574 60004 54626
rect 59948 54292 60004 54574
rect 59948 54226 60004 54236
rect 60060 54514 60116 54526
rect 60060 54462 60062 54514
rect 60114 54462 60116 54514
rect 60060 53954 60116 54462
rect 60060 53902 60062 53954
rect 60114 53902 60116 53954
rect 60060 53890 60116 53902
rect 60172 51602 60228 61068
rect 60396 61058 60452 61068
rect 60396 60676 60452 60686
rect 60284 59106 60340 59118
rect 60284 59054 60286 59106
rect 60338 59054 60340 59106
rect 60284 58434 60340 59054
rect 60284 58382 60286 58434
rect 60338 58382 60340 58434
rect 60284 58370 60340 58382
rect 60396 57988 60452 60620
rect 60508 59892 60564 63870
rect 61180 63924 61236 63934
rect 61180 63830 61236 63868
rect 61740 61684 61796 64204
rect 61964 63252 62020 64204
rect 61852 63196 62020 63252
rect 61852 62580 61908 63196
rect 62412 63138 62468 63150
rect 62412 63086 62414 63138
rect 62466 63086 62468 63138
rect 61964 63028 62020 63038
rect 61964 63026 62132 63028
rect 61964 62974 61966 63026
rect 62018 62974 62132 63026
rect 61964 62972 62132 62974
rect 61964 62962 62020 62972
rect 61964 62580 62020 62590
rect 61852 62578 62020 62580
rect 61852 62526 61966 62578
rect 62018 62526 62020 62578
rect 61852 62524 62020 62526
rect 61964 62514 62020 62524
rect 61852 62354 61908 62366
rect 61852 62302 61854 62354
rect 61906 62302 61908 62354
rect 61852 61908 61908 62302
rect 62076 61908 62132 62972
rect 62300 63026 62356 63038
rect 62300 62974 62302 63026
rect 62354 62974 62356 63026
rect 62188 62916 62244 62926
rect 62188 62822 62244 62860
rect 62188 62468 62244 62478
rect 62300 62468 62356 62974
rect 62244 62412 62356 62468
rect 62412 62468 62468 63086
rect 62972 62916 63028 62926
rect 62972 62914 63140 62916
rect 62972 62862 62974 62914
rect 63026 62862 63140 62914
rect 62972 62860 63140 62862
rect 62972 62850 63028 62860
rect 62972 62468 63028 62478
rect 62412 62466 63028 62468
rect 62412 62414 62414 62466
rect 62466 62414 62974 62466
rect 63026 62414 63028 62466
rect 62412 62412 63028 62414
rect 63084 62468 63140 62860
rect 63420 62914 63476 62926
rect 63420 62862 63422 62914
rect 63474 62862 63476 62914
rect 63308 62580 63364 62590
rect 63308 62486 63364 62524
rect 63196 62468 63252 62478
rect 63084 62412 63196 62468
rect 62188 62374 62244 62412
rect 62412 62402 62468 62412
rect 62860 61908 62916 61918
rect 62076 61852 62468 61908
rect 61852 61842 61908 61852
rect 61740 61628 62020 61684
rect 61852 61460 61908 61470
rect 61740 61458 61908 61460
rect 61740 61406 61854 61458
rect 61906 61406 61908 61458
rect 61740 61404 61908 61406
rect 61628 61348 61684 61358
rect 60508 59826 60564 59836
rect 61404 60674 61460 60686
rect 61404 60622 61406 60674
rect 61458 60622 61460 60674
rect 61068 59444 61124 59454
rect 60956 58436 61012 58446
rect 60620 58324 60676 58334
rect 60620 58230 60676 58268
rect 60284 57932 60452 57988
rect 60508 58210 60564 58222
rect 60508 58158 60510 58210
rect 60562 58158 60564 58210
rect 60284 55468 60340 57932
rect 60396 57650 60452 57662
rect 60396 57598 60398 57650
rect 60450 57598 60452 57650
rect 60396 57092 60452 57598
rect 60396 57026 60452 57036
rect 60284 55412 60452 55468
rect 60284 53954 60340 53966
rect 60284 53902 60286 53954
rect 60338 53902 60340 53954
rect 60284 53506 60340 53902
rect 60284 53454 60286 53506
rect 60338 53454 60340 53506
rect 60284 52948 60340 53454
rect 60284 52882 60340 52892
rect 60172 51550 60174 51602
rect 60226 51550 60228 51602
rect 60172 51538 60228 51550
rect 59724 51492 59780 51502
rect 59724 51398 59780 51436
rect 60284 51380 60340 51390
rect 60284 51286 60340 51324
rect 59724 50820 59780 50830
rect 59724 50706 59780 50764
rect 59724 50654 59726 50706
rect 59778 50654 59780 50706
rect 59724 50642 59780 50654
rect 60172 50708 60228 50718
rect 60172 50614 60228 50652
rect 59724 48132 59780 48142
rect 59724 48038 59780 48076
rect 59948 47572 60004 47582
rect 59948 47478 60004 47516
rect 59612 43810 59668 43820
rect 59836 43652 59892 43662
rect 58492 43598 58494 43650
rect 58546 43598 58548 43650
rect 58492 43586 58548 43598
rect 59612 43650 59892 43652
rect 59612 43598 59838 43650
rect 59890 43598 59892 43650
rect 59612 43596 59892 43598
rect 58716 43538 58772 43550
rect 58716 43486 58718 43538
rect 58770 43486 58772 43538
rect 58716 43428 58772 43486
rect 58716 43362 58772 43372
rect 59276 43428 59332 43438
rect 59276 43334 59332 43372
rect 58940 42868 58996 42878
rect 58940 41410 58996 42812
rect 58940 41358 58942 41410
rect 58994 41358 58996 41410
rect 58940 41346 58996 41358
rect 58604 41188 58660 41198
rect 58604 41094 58660 41132
rect 59500 41074 59556 41086
rect 59500 41022 59502 41074
rect 59554 41022 59556 41074
rect 59500 40964 59556 41022
rect 59500 40898 59556 40908
rect 59612 40514 59668 43596
rect 59836 43586 59892 43596
rect 60172 43538 60228 43550
rect 60172 43486 60174 43538
rect 60226 43486 60228 43538
rect 60172 41860 60228 43486
rect 60396 43316 60452 55412
rect 60508 55076 60564 58158
rect 60956 57764 61012 58380
rect 60732 57762 61012 57764
rect 60732 57710 60958 57762
rect 61010 57710 61012 57762
rect 60732 57708 61012 57710
rect 60620 57092 60676 57102
rect 60620 55524 60676 57036
rect 60620 55298 60676 55468
rect 60620 55246 60622 55298
rect 60674 55246 60676 55298
rect 60620 55234 60676 55246
rect 60508 55010 60564 55020
rect 60732 54514 60788 57708
rect 60956 57698 61012 57708
rect 61068 56644 61124 59388
rect 61404 58546 61460 60622
rect 61628 59220 61684 61292
rect 61740 60564 61796 61404
rect 61852 61394 61908 61404
rect 61852 60900 61908 60910
rect 61852 60786 61908 60844
rect 61852 60734 61854 60786
rect 61906 60734 61908 60786
rect 61852 60722 61908 60734
rect 61964 60788 62020 61628
rect 62300 61570 62356 61582
rect 62300 61518 62302 61570
rect 62354 61518 62356 61570
rect 62300 60900 62356 61518
rect 62412 61010 62468 61852
rect 62748 61684 62804 61694
rect 62748 61570 62804 61628
rect 62748 61518 62750 61570
rect 62802 61518 62804 61570
rect 62748 61506 62804 61518
rect 62860 61458 62916 61852
rect 62972 61572 63028 62412
rect 63196 62374 63252 62412
rect 63420 62468 63476 62862
rect 63420 62402 63476 62412
rect 62972 61506 63028 61516
rect 63532 62354 63588 62366
rect 63532 62302 63534 62354
rect 63586 62302 63588 62354
rect 62860 61406 62862 61458
rect 62914 61406 62916 61458
rect 62860 61394 62916 61406
rect 63308 61458 63364 61470
rect 63308 61406 63310 61458
rect 63362 61406 63364 61458
rect 62412 60958 62414 61010
rect 62466 60958 62468 61010
rect 62412 60946 62468 60958
rect 62300 60834 62356 60844
rect 62188 60788 62244 60798
rect 61964 60786 62244 60788
rect 61964 60734 62190 60786
rect 62242 60734 62244 60786
rect 61964 60732 62244 60734
rect 62188 60722 62244 60732
rect 63084 60788 63140 60798
rect 63308 60788 63364 61406
rect 63084 60786 63364 60788
rect 63084 60734 63086 60786
rect 63138 60734 63364 60786
rect 63084 60732 63364 60734
rect 61740 60508 61908 60564
rect 61740 59778 61796 59790
rect 61740 59726 61742 59778
rect 61794 59726 61796 59778
rect 61740 59444 61796 59726
rect 61740 59378 61796 59388
rect 61628 59164 61796 59220
rect 61404 58494 61406 58546
rect 61458 58494 61460 58546
rect 61404 57876 61460 58494
rect 61404 57810 61460 57820
rect 60732 54462 60734 54514
rect 60786 54462 60788 54514
rect 60732 54450 60788 54462
rect 60844 56588 61124 56644
rect 61516 56866 61572 56878
rect 61516 56814 61518 56866
rect 61570 56814 61572 56866
rect 60844 56194 60900 56588
rect 60844 56142 60846 56194
rect 60898 56142 60900 56194
rect 60844 55188 60900 56142
rect 60956 56196 61012 56206
rect 60956 56194 61460 56196
rect 60956 56142 60958 56194
rect 61010 56142 61460 56194
rect 60956 56140 61460 56142
rect 60956 56130 61012 56140
rect 60844 53172 60900 55132
rect 60956 55858 61012 55870
rect 60956 55806 60958 55858
rect 61010 55806 61012 55858
rect 60956 53844 61012 55806
rect 61180 55412 61236 55422
rect 60956 53778 61012 53788
rect 61068 54516 61124 54526
rect 60844 53106 60900 53116
rect 61068 52836 61124 54460
rect 61180 53060 61236 55356
rect 61292 55188 61348 55198
rect 61292 55094 61348 55132
rect 61404 54852 61460 56140
rect 61292 54796 61460 54852
rect 61516 56084 61572 56814
rect 61628 56084 61684 56094
rect 61516 56082 61684 56084
rect 61516 56030 61630 56082
rect 61682 56030 61684 56082
rect 61516 56028 61684 56030
rect 61516 55188 61572 56028
rect 61628 56018 61684 56028
rect 61292 53508 61348 54796
rect 61404 54628 61460 54638
rect 61404 54534 61460 54572
rect 61516 53730 61572 55132
rect 61516 53678 61518 53730
rect 61570 53678 61572 53730
rect 61516 53666 61572 53678
rect 61292 53452 61684 53508
rect 61628 53170 61684 53452
rect 61628 53118 61630 53170
rect 61682 53118 61684 53170
rect 61628 53106 61684 53118
rect 61180 53004 61460 53060
rect 61180 52836 61236 52846
rect 60508 52834 61236 52836
rect 60508 52782 61182 52834
rect 61234 52782 61236 52834
rect 60508 52780 61236 52782
rect 60508 47572 60564 52780
rect 61180 52770 61236 52780
rect 60844 51940 60900 51950
rect 60844 51380 60900 51884
rect 60844 51286 60900 51324
rect 61180 51268 61236 51278
rect 60620 48804 60676 48814
rect 60620 48710 60676 48748
rect 60732 48356 60788 48366
rect 60732 48354 60900 48356
rect 60732 48302 60734 48354
rect 60786 48302 60900 48354
rect 60732 48300 60900 48302
rect 60732 48290 60788 48300
rect 60620 48244 60676 48254
rect 60620 48150 60676 48188
rect 60844 48020 60900 48300
rect 60844 47954 60900 47964
rect 60956 48242 61012 48254
rect 60956 48190 60958 48242
rect 61010 48190 61012 48242
rect 60620 47572 60676 47582
rect 60508 47570 60676 47572
rect 60508 47518 60622 47570
rect 60674 47518 60676 47570
rect 60508 47516 60676 47518
rect 60620 47460 60676 47516
rect 60620 47394 60676 47404
rect 60956 46788 61012 48190
rect 60956 46722 61012 46732
rect 61068 47348 61124 47358
rect 60956 46564 61012 46574
rect 61068 46564 61124 47292
rect 60956 46562 61124 46564
rect 60956 46510 60958 46562
rect 61010 46510 61124 46562
rect 60956 46508 61124 46510
rect 60956 46498 61012 46508
rect 60396 43250 60452 43260
rect 60396 42868 60452 42878
rect 60396 42774 60452 42812
rect 60172 41794 60228 41804
rect 60732 42082 60788 42094
rect 60732 42030 60734 42082
rect 60786 42030 60788 42082
rect 60732 41972 60788 42030
rect 59724 41188 59780 41198
rect 60284 41188 60340 41198
rect 59724 41186 60340 41188
rect 59724 41134 59726 41186
rect 59778 41134 60286 41186
rect 60338 41134 60340 41186
rect 59724 41132 60340 41134
rect 59724 41122 59780 41132
rect 59612 40462 59614 40514
rect 59666 40462 59668 40514
rect 59612 40450 59668 40462
rect 58940 40404 58996 40414
rect 58716 40348 58940 40404
rect 58716 38834 58772 40348
rect 58940 40310 58996 40348
rect 59948 39506 60004 39518
rect 59948 39454 59950 39506
rect 60002 39454 60004 39506
rect 59612 39396 59668 39406
rect 59388 39394 59668 39396
rect 59388 39342 59614 39394
rect 59666 39342 59668 39394
rect 59388 39340 59668 39342
rect 59388 38946 59444 39340
rect 59612 39330 59668 39340
rect 59948 39060 60004 39454
rect 60284 39396 60340 41132
rect 60732 39620 60788 41916
rect 60732 39554 60788 39564
rect 60284 39330 60340 39340
rect 59948 38994 60004 39004
rect 59388 38894 59390 38946
rect 59442 38894 59444 38946
rect 59388 38882 59444 38894
rect 58716 38782 58718 38834
rect 58770 38782 58772 38834
rect 58716 38770 58772 38782
rect 61068 38164 61124 38174
rect 58716 37716 58772 37726
rect 58716 37268 58772 37660
rect 59388 37716 59444 37726
rect 58828 37492 58884 37502
rect 58828 37380 58884 37436
rect 59388 37490 59444 37660
rect 59388 37438 59390 37490
rect 59442 37438 59444 37490
rect 59388 37426 59444 37438
rect 59724 37716 59780 37726
rect 58828 37378 58996 37380
rect 58828 37326 58830 37378
rect 58882 37326 58996 37378
rect 58828 37324 58996 37326
rect 58828 37314 58884 37324
rect 58492 37266 58772 37268
rect 58492 37214 58718 37266
rect 58770 37214 58772 37266
rect 58492 37212 58772 37214
rect 58492 35810 58548 37212
rect 58716 37202 58772 37212
rect 58940 36594 58996 37324
rect 58940 36542 58942 36594
rect 58994 36542 58996 36594
rect 58940 36530 58996 36542
rect 59500 36372 59556 36382
rect 59052 36370 59556 36372
rect 59052 36318 59502 36370
rect 59554 36318 59556 36370
rect 59052 36316 59556 36318
rect 59052 35922 59108 36316
rect 59500 36306 59556 36316
rect 59052 35870 59054 35922
rect 59106 35870 59108 35922
rect 59052 35858 59108 35870
rect 59724 35922 59780 37660
rect 59836 37492 59892 37502
rect 59836 37398 59892 37436
rect 59724 35870 59726 35922
rect 59778 35870 59780 35922
rect 59724 35858 59780 35870
rect 59836 36258 59892 36270
rect 59836 36206 59838 36258
rect 59890 36206 59892 36258
rect 58492 35758 58494 35810
rect 58546 35758 58548 35810
rect 58492 35746 58548 35758
rect 58604 35812 58660 35822
rect 58380 33954 58436 33964
rect 58604 33572 58660 35756
rect 58716 35476 58772 35486
rect 58716 35382 58772 35420
rect 59612 34244 59668 34254
rect 59836 34244 59892 36206
rect 60284 36260 60340 36270
rect 60284 36258 60452 36260
rect 60284 36206 60286 36258
rect 60338 36206 60452 36258
rect 60284 36204 60452 36206
rect 60284 36194 60340 36204
rect 60284 35700 60340 35710
rect 60284 35606 60340 35644
rect 59612 34242 59892 34244
rect 59612 34190 59614 34242
rect 59666 34190 59892 34242
rect 59612 34188 59892 34190
rect 59948 34692 60004 34702
rect 59612 34178 59668 34188
rect 58604 33516 58996 33572
rect 58380 33348 58436 33358
rect 58380 33254 58436 33292
rect 58940 33234 58996 33516
rect 59724 33460 59780 33470
rect 59948 33460 60004 34636
rect 60284 34132 60340 34142
rect 60396 34132 60452 36204
rect 61068 35922 61124 38108
rect 61180 37492 61236 51212
rect 61292 49698 61348 49710
rect 61292 49646 61294 49698
rect 61346 49646 61348 49698
rect 61292 47348 61348 49646
rect 61404 49138 61460 53004
rect 61628 52276 61684 52286
rect 61628 51602 61684 52220
rect 61628 51550 61630 51602
rect 61682 51550 61684 51602
rect 61628 51380 61684 51550
rect 61628 51314 61684 51324
rect 61740 51156 61796 59164
rect 61852 59108 61908 60508
rect 62860 60002 62916 60014
rect 62860 59950 62862 60002
rect 62914 59950 62916 60002
rect 62188 59780 62244 59790
rect 62860 59780 62916 59950
rect 63084 60004 63140 60732
rect 63532 60564 63588 62302
rect 63644 61348 63700 68796
rect 63756 68292 63812 71596
rect 65324 71652 65380 72156
rect 65324 71586 65380 71596
rect 65436 72324 65492 72334
rect 64316 71092 64372 71102
rect 64316 70998 64372 71036
rect 64764 70754 64820 70766
rect 65324 70756 65380 70766
rect 64764 70702 64766 70754
rect 64818 70702 64820 70754
rect 63868 70420 63924 70430
rect 63868 69522 63924 70364
rect 64764 70420 64820 70702
rect 64764 70354 64820 70364
rect 64876 70754 65380 70756
rect 64876 70702 65326 70754
rect 65378 70702 65380 70754
rect 64876 70700 65380 70702
rect 63868 69470 63870 69522
rect 63922 69470 63924 69522
rect 63868 69458 63924 69470
rect 63868 68628 63924 68638
rect 63868 68534 63924 68572
rect 64316 68514 64372 68526
rect 64316 68462 64318 68514
rect 64370 68462 64372 68514
rect 63756 68236 63924 68292
rect 63756 68068 63812 68078
rect 63756 61684 63812 68012
rect 63868 61796 63924 68236
rect 64316 68068 64372 68462
rect 64316 68002 64372 68012
rect 64876 67954 64932 70700
rect 65324 70690 65380 70700
rect 65436 70532 65492 72268
rect 64876 67902 64878 67954
rect 64930 67902 64932 67954
rect 64876 67890 64932 67902
rect 65212 70476 65492 70532
rect 64092 67842 64148 67854
rect 64092 67790 64094 67842
rect 64146 67790 64148 67842
rect 64092 64708 64148 67790
rect 64988 66050 65044 66062
rect 64988 65998 64990 66050
rect 65042 65998 65044 66050
rect 64988 65716 65044 65998
rect 64988 65650 65044 65660
rect 64316 65604 64372 65614
rect 64316 65510 64372 65548
rect 64652 65602 64708 65614
rect 64652 65550 64654 65602
rect 64706 65550 64708 65602
rect 64652 64820 64708 65550
rect 64764 64820 64820 64830
rect 64652 64818 64820 64820
rect 64652 64766 64766 64818
rect 64818 64766 64820 64818
rect 64652 64764 64820 64766
rect 64764 64754 64820 64764
rect 64092 64614 64148 64652
rect 63980 62580 64036 62590
rect 63980 62486 64036 62524
rect 64876 62244 64932 62254
rect 65212 62188 65268 70476
rect 63868 61740 64036 61796
rect 63756 61618 63812 61628
rect 63644 61292 63812 61348
rect 63644 61124 63700 61134
rect 63644 60786 63700 61068
rect 63644 60734 63646 60786
rect 63698 60734 63700 60786
rect 63644 60722 63700 60734
rect 63532 60498 63588 60508
rect 63644 60116 63700 60126
rect 63644 60004 63700 60060
rect 63084 59938 63140 59948
rect 63532 60002 63700 60004
rect 63532 59950 63646 60002
rect 63698 59950 63700 60002
rect 63532 59948 63700 59950
rect 62188 59778 62916 59780
rect 62188 59726 62190 59778
rect 62242 59726 62916 59778
rect 62188 59724 62916 59726
rect 62188 59714 62244 59724
rect 62860 59556 62916 59724
rect 62860 59500 63364 59556
rect 63084 59332 63140 59342
rect 62972 59330 63140 59332
rect 62972 59278 63086 59330
rect 63138 59278 63140 59330
rect 62972 59276 63140 59278
rect 62860 59220 62916 59230
rect 62524 59218 62916 59220
rect 62524 59166 62862 59218
rect 62914 59166 62916 59218
rect 62524 59164 62916 59166
rect 61852 59042 61908 59052
rect 62412 59108 62468 59118
rect 62412 59014 62468 59052
rect 62524 57988 62580 59164
rect 62860 59154 62916 59164
rect 62188 57932 62580 57988
rect 62748 58996 62804 59006
rect 62188 56978 62244 57932
rect 62188 56926 62190 56978
rect 62242 56926 62244 56978
rect 62188 56914 62244 56926
rect 62412 55970 62468 55982
rect 62412 55918 62414 55970
rect 62466 55918 62468 55970
rect 62412 55412 62468 55918
rect 62412 55346 62468 55356
rect 62412 55186 62468 55198
rect 62412 55134 62414 55186
rect 62466 55134 62468 55186
rect 62076 55074 62132 55086
rect 62076 55022 62078 55074
rect 62130 55022 62132 55074
rect 62076 54628 62132 55022
rect 62300 55074 62356 55086
rect 62300 55022 62302 55074
rect 62354 55022 62356 55074
rect 62300 54740 62356 55022
rect 62412 55076 62468 55134
rect 62412 55010 62468 55020
rect 62300 54674 62356 54684
rect 62076 54562 62132 54572
rect 61852 54516 61908 54526
rect 61852 53170 61908 54460
rect 62188 53844 62244 53854
rect 62188 53730 62244 53788
rect 62188 53678 62190 53730
rect 62242 53678 62244 53730
rect 62188 53666 62244 53678
rect 61852 53118 61854 53170
rect 61906 53118 61908 53170
rect 61852 53106 61908 53118
rect 62636 53058 62692 53070
rect 62636 53006 62638 53058
rect 62690 53006 62692 53058
rect 61964 52948 62020 52958
rect 61964 52854 62020 52892
rect 62524 52948 62580 52958
rect 62076 52388 62132 52398
rect 62076 51602 62132 52332
rect 62076 51550 62078 51602
rect 62130 51550 62132 51602
rect 62076 51492 62132 51550
rect 62076 51426 62132 51436
rect 62188 52386 62244 52398
rect 62188 52334 62190 52386
rect 62242 52334 62244 52386
rect 62188 52274 62244 52334
rect 62188 52222 62190 52274
rect 62242 52222 62244 52274
rect 61740 51090 61796 51100
rect 61404 49086 61406 49138
rect 61458 49086 61460 49138
rect 61404 47572 61460 49086
rect 61852 50594 61908 50606
rect 61852 50542 61854 50594
rect 61906 50542 61908 50594
rect 61852 49810 61908 50542
rect 61852 49758 61854 49810
rect 61906 49758 61908 49810
rect 61852 48916 61908 49758
rect 61404 47506 61460 47516
rect 61628 48860 61852 48916
rect 61516 47460 61572 47470
rect 61404 47348 61460 47358
rect 61292 47292 61404 47348
rect 61404 47254 61460 47292
rect 61516 47346 61572 47404
rect 61516 47294 61518 47346
rect 61570 47294 61572 47346
rect 61516 47282 61572 47294
rect 61516 46676 61572 46686
rect 61628 46676 61684 48860
rect 61852 48850 61908 48860
rect 61964 49924 62020 49934
rect 61740 48468 61796 48478
rect 61740 47458 61796 48412
rect 61852 48468 61908 48478
rect 61964 48468 62020 49868
rect 62188 48804 62244 52222
rect 62524 52164 62580 52892
rect 62636 52386 62692 53006
rect 62636 52334 62638 52386
rect 62690 52334 62692 52386
rect 62636 52322 62692 52334
rect 62636 52164 62692 52174
rect 62524 52108 62636 52164
rect 62636 52070 62692 52108
rect 62636 51268 62692 51278
rect 62188 48738 62244 48748
rect 62412 51266 62692 51268
rect 62412 51214 62638 51266
rect 62690 51214 62692 51266
rect 62412 51212 62692 51214
rect 62412 51044 62468 51212
rect 62636 51202 62692 51212
rect 61852 48466 62132 48468
rect 61852 48414 61854 48466
rect 61906 48414 62132 48466
rect 61852 48412 62132 48414
rect 61852 48402 61908 48412
rect 61964 48242 62020 48254
rect 61964 48190 61966 48242
rect 62018 48190 62020 48242
rect 61852 48020 61908 48030
rect 61852 47926 61908 47964
rect 61740 47406 61742 47458
rect 61794 47406 61796 47458
rect 61740 47394 61796 47406
rect 61852 47572 61908 47582
rect 61516 46674 61684 46676
rect 61516 46622 61518 46674
rect 61570 46622 61684 46674
rect 61516 46620 61684 46622
rect 61516 45890 61572 46620
rect 61516 45838 61518 45890
rect 61570 45838 61572 45890
rect 61516 45826 61572 45838
rect 61404 44996 61460 45006
rect 61404 44902 61460 44940
rect 61852 44434 61908 47516
rect 61964 47348 62020 48190
rect 62076 47570 62132 48412
rect 62076 47518 62078 47570
rect 62130 47518 62132 47570
rect 62076 47506 62132 47518
rect 62300 48020 62356 48030
rect 61964 47282 62020 47292
rect 62188 46788 62244 46798
rect 62188 46694 62244 46732
rect 62188 46004 62244 46014
rect 62300 46004 62356 47964
rect 62188 46002 62356 46004
rect 62188 45950 62190 46002
rect 62242 45950 62356 46002
rect 62188 45948 62356 45950
rect 62188 45938 62244 45948
rect 61852 44382 61854 44434
rect 61906 44382 61908 44434
rect 61852 44212 61908 44382
rect 61292 42530 61348 42542
rect 61292 42478 61294 42530
rect 61346 42478 61348 42530
rect 61292 41972 61348 42478
rect 61292 41906 61348 41916
rect 61852 41972 61908 44156
rect 61852 41906 61908 41916
rect 62076 43316 62132 43326
rect 62076 42530 62132 43260
rect 62076 42478 62078 42530
rect 62130 42478 62132 42530
rect 62076 41970 62132 42478
rect 62076 41918 62078 41970
rect 62130 41918 62132 41970
rect 62076 41906 62132 41918
rect 62412 42868 62468 50988
rect 62636 50484 62692 50494
rect 62636 50390 62692 50428
rect 62524 49812 62580 49822
rect 62524 49718 62580 49756
rect 62636 48804 62692 48814
rect 62524 48580 62580 48590
rect 62524 48354 62580 48524
rect 62636 48466 62692 48748
rect 62636 48414 62638 48466
rect 62690 48414 62692 48466
rect 62636 48402 62692 48414
rect 62748 48692 62804 58940
rect 62972 55468 63028 59276
rect 63084 59266 63140 59276
rect 63196 59218 63252 59230
rect 63196 59166 63198 59218
rect 63250 59166 63252 59218
rect 63196 58660 63252 59166
rect 63196 58594 63252 58604
rect 62972 55412 63140 55468
rect 63084 54740 63140 55412
rect 63084 54674 63140 54684
rect 62860 54628 62916 54638
rect 62860 53170 62916 54572
rect 62860 53118 62862 53170
rect 62914 53118 62916 53170
rect 62860 53106 62916 53118
rect 63196 53172 63252 53182
rect 63196 53078 63252 53116
rect 62972 51268 63028 51278
rect 62972 51174 63028 51212
rect 62524 48302 62526 48354
rect 62578 48302 62580 48354
rect 62524 47348 62580 48302
rect 62748 47572 62804 48636
rect 63196 50484 63252 50494
rect 63196 48466 63252 50428
rect 63196 48414 63198 48466
rect 63250 48414 63252 48466
rect 63196 48402 63252 48414
rect 62860 48356 62916 48366
rect 62860 48262 62916 48300
rect 62860 47572 62916 47582
rect 62748 47570 62916 47572
rect 62748 47518 62862 47570
rect 62914 47518 62916 47570
rect 62748 47516 62916 47518
rect 62860 47506 62916 47516
rect 62524 47282 62580 47292
rect 62524 44322 62580 44334
rect 62524 44270 62526 44322
rect 62578 44270 62580 44322
rect 62524 43764 62580 44270
rect 62524 43698 62580 43708
rect 62748 44098 62804 44110
rect 62748 44046 62750 44098
rect 62802 44046 62804 44098
rect 62524 42868 62580 42878
rect 62412 42866 62580 42868
rect 62412 42814 62526 42866
rect 62578 42814 62580 42866
rect 62412 42812 62580 42814
rect 61740 41748 61796 41758
rect 61292 40404 61348 40414
rect 61292 39394 61348 40348
rect 61740 40290 61796 41692
rect 62412 41748 62468 42812
rect 62524 42802 62580 42812
rect 62748 42868 62804 44046
rect 62748 42802 62804 42812
rect 62412 41682 62468 41692
rect 63084 42754 63140 42766
rect 63084 42702 63086 42754
rect 63138 42702 63140 42754
rect 62188 41300 62244 41310
rect 62188 41206 62244 41244
rect 63084 41188 63140 42702
rect 62748 41076 62804 41086
rect 62188 40628 62244 40638
rect 62188 40534 62244 40572
rect 62748 40626 62804 41020
rect 62748 40574 62750 40626
rect 62802 40574 62804 40626
rect 62748 40516 62804 40574
rect 63084 40628 63140 41132
rect 63084 40562 63140 40572
rect 62748 40450 62804 40460
rect 61740 40238 61742 40290
rect 61794 40238 61796 40290
rect 61740 40226 61796 40238
rect 61292 39342 61294 39394
rect 61346 39342 61348 39394
rect 61292 38052 61348 39342
rect 61740 39620 61796 39630
rect 61516 38724 61572 38734
rect 61516 38630 61572 38668
rect 61516 38164 61572 38174
rect 61516 38070 61572 38108
rect 61348 37996 61460 38052
rect 61292 37986 61348 37996
rect 61180 37426 61236 37436
rect 61068 35870 61070 35922
rect 61122 35870 61124 35922
rect 60620 35810 60676 35822
rect 60620 35758 60622 35810
rect 60674 35758 60676 35810
rect 60620 35028 60676 35758
rect 61068 35812 61124 35870
rect 61068 35746 61124 35756
rect 60620 34962 60676 34972
rect 61404 34914 61460 37996
rect 61516 37828 61572 37838
rect 61516 37044 61572 37772
rect 61516 36594 61572 36988
rect 61516 36542 61518 36594
rect 61570 36542 61572 36594
rect 61516 36530 61572 36542
rect 61740 35588 61796 39564
rect 62300 39620 62356 39630
rect 62300 39526 62356 39564
rect 62524 39396 62580 39406
rect 62188 39060 62244 39070
rect 62188 38966 62244 39004
rect 62524 38834 62580 39340
rect 63196 39284 63252 39294
rect 62524 38782 62526 38834
rect 62578 38782 62580 38834
rect 62524 38724 62580 38782
rect 62524 38658 62580 38668
rect 62860 38948 62916 38958
rect 62860 38162 62916 38892
rect 62860 38110 62862 38162
rect 62914 38110 62916 38162
rect 62860 38098 62916 38110
rect 63084 38946 63140 38958
rect 63084 38894 63086 38946
rect 63138 38894 63140 38946
rect 63084 38164 63140 38894
rect 63196 38834 63252 39228
rect 63196 38782 63198 38834
rect 63250 38782 63252 38834
rect 63196 38724 63252 38782
rect 63196 38658 63252 38668
rect 63084 38098 63140 38108
rect 62188 38052 62244 38062
rect 62188 37958 62244 37996
rect 61964 37044 62020 37054
rect 61964 35810 62020 36988
rect 62748 36036 62804 36046
rect 61964 35758 61966 35810
rect 62018 35758 62020 35810
rect 61964 35746 62020 35758
rect 62524 35810 62580 35822
rect 62524 35758 62526 35810
rect 62578 35758 62580 35810
rect 61404 34862 61406 34914
rect 61458 34862 61460 34914
rect 61404 34850 61460 34862
rect 61516 35532 61740 35588
rect 60340 34076 60452 34132
rect 60732 34132 60788 34142
rect 60284 34038 60340 34076
rect 59724 33458 60004 33460
rect 59724 33406 59726 33458
rect 59778 33406 60004 33458
rect 59724 33404 60004 33406
rect 59164 33348 59220 33358
rect 59164 33254 59220 33292
rect 59724 33348 59780 33404
rect 59724 33282 59780 33292
rect 60396 33346 60452 33358
rect 60396 33294 60398 33346
rect 60450 33294 60452 33346
rect 58940 33182 58942 33234
rect 58994 33182 58996 33234
rect 58380 32788 58436 32798
rect 58268 32786 58436 32788
rect 58268 32734 58382 32786
rect 58434 32734 58436 32786
rect 58268 32732 58436 32734
rect 58380 32722 58436 32732
rect 58940 32788 58996 33182
rect 58940 32722 58996 32732
rect 59724 32788 59780 32798
rect 59724 32694 59780 32732
rect 60396 32788 60452 33294
rect 60620 33236 60676 33246
rect 60620 33142 60676 33180
rect 60396 32722 60452 32732
rect 60732 32788 60788 34076
rect 60956 34132 61012 34142
rect 60956 34038 61012 34076
rect 61404 33460 61460 33470
rect 61516 33460 61572 35532
rect 61740 35522 61796 35532
rect 62188 35028 62244 35038
rect 62188 34934 62244 34972
rect 62524 35028 62580 35758
rect 62748 35698 62804 35980
rect 62748 35646 62750 35698
rect 62802 35646 62804 35698
rect 62748 35634 62804 35646
rect 63084 35700 63140 35710
rect 63084 35606 63140 35644
rect 62524 34962 62580 34972
rect 62188 34356 62244 34366
rect 61404 33458 61572 33460
rect 61404 33406 61406 33458
rect 61458 33406 61572 33458
rect 61404 33404 61572 33406
rect 61740 34018 61796 34030
rect 61740 33966 61742 34018
rect 61794 33966 61796 34018
rect 61404 33394 61460 33404
rect 61740 33236 61796 33966
rect 61740 33170 61796 33180
rect 61964 34020 62020 34030
rect 61068 32788 61124 32798
rect 60732 32786 61124 32788
rect 60732 32734 60734 32786
rect 60786 32734 61070 32786
rect 61122 32734 61124 32786
rect 60732 32732 61124 32734
rect 60732 32722 60788 32732
rect 61068 32722 61124 32732
rect 61740 32788 61796 32798
rect 61740 32694 61796 32732
rect 57932 31838 57934 31890
rect 57986 31838 57988 31890
rect 57932 31826 57988 31838
rect 61404 32676 61460 32686
rect 61404 31890 61460 32620
rect 61964 32564 62020 33964
rect 62188 33684 62244 34300
rect 63308 34356 63364 59500
rect 63532 58996 63588 59948
rect 63644 59938 63700 59948
rect 63532 58930 63588 58940
rect 63644 59218 63700 59230
rect 63644 59166 63646 59218
rect 63698 59166 63700 59218
rect 63532 58548 63588 58558
rect 63644 58548 63700 59166
rect 63532 58546 63700 58548
rect 63532 58494 63534 58546
rect 63586 58494 63700 58546
rect 63532 58492 63700 58494
rect 63532 58482 63588 58492
rect 63532 56196 63588 56206
rect 63532 54402 63588 56140
rect 63532 54350 63534 54402
rect 63586 54350 63588 54402
rect 63532 54338 63588 54350
rect 63420 53172 63476 53182
rect 63420 53078 63476 53116
rect 63532 53060 63588 53070
rect 63532 52966 63588 53004
rect 63756 51940 63812 61292
rect 63980 60676 64036 61740
rect 63980 60610 64036 60620
rect 64092 61570 64148 61582
rect 64876 61572 64932 62188
rect 64092 61518 64094 61570
rect 64146 61518 64148 61570
rect 64092 61012 64148 61518
rect 63868 59444 63924 59454
rect 63868 59350 63924 59388
rect 63980 59220 64036 59230
rect 63980 59126 64036 59164
rect 63980 55412 64036 55422
rect 63868 55188 63924 55198
rect 63868 55094 63924 55132
rect 63980 54738 64036 55356
rect 63980 54686 63982 54738
rect 64034 54686 64036 54738
rect 63980 54674 64036 54686
rect 63980 52834 64036 52846
rect 63980 52782 63982 52834
rect 64034 52782 64036 52834
rect 63980 52164 64036 52782
rect 63980 52098 64036 52108
rect 63756 51874 63812 51884
rect 63980 51604 64036 51614
rect 64092 51604 64148 60956
rect 64764 61570 64932 61572
rect 64764 61518 64878 61570
rect 64930 61518 64932 61570
rect 64764 61516 64932 61518
rect 64540 60788 64596 60798
rect 64540 60694 64596 60732
rect 64428 60004 64484 60014
rect 64428 59910 64484 59948
rect 64764 59780 64820 61516
rect 64876 61506 64932 61516
rect 65100 62132 65268 62188
rect 65324 70308 65380 70318
rect 65324 62188 65380 70252
rect 65436 69412 65492 69422
rect 65436 68964 65492 69356
rect 65436 65716 65492 68908
rect 65548 68852 65604 73500
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 65772 72324 65828 72334
rect 65772 72230 65828 72268
rect 66108 71650 66164 71662
rect 66108 71598 66110 71650
rect 66162 71598 66164 71650
rect 66108 71540 66164 71598
rect 66108 71484 66388 71540
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 65660 70868 65716 70878
rect 65660 70866 66276 70868
rect 65660 70814 65662 70866
rect 65714 70814 66276 70866
rect 65660 70812 66276 70814
rect 65660 70802 65716 70812
rect 66220 70418 66276 70812
rect 66332 70866 66388 71484
rect 67228 71092 67284 75964
rect 67340 75908 67396 76414
rect 67340 75842 67396 75852
rect 66332 70814 66334 70866
rect 66386 70814 66388 70866
rect 66332 70756 66388 70814
rect 66668 71090 67396 71092
rect 66668 71038 67230 71090
rect 67282 71038 67396 71090
rect 66668 71036 67396 71038
rect 66668 70866 66724 71036
rect 67228 71026 67284 71036
rect 66668 70814 66670 70866
rect 66722 70814 66724 70866
rect 66668 70802 66724 70814
rect 66332 70690 66388 70700
rect 66220 70366 66222 70418
rect 66274 70366 66276 70418
rect 66220 70354 66276 70366
rect 66780 70308 66836 70318
rect 66780 70214 66836 70252
rect 67340 70308 67396 71036
rect 67452 70532 67508 79662
rect 68124 79602 68180 81004
rect 68236 80164 68292 81676
rect 68348 81730 68404 81742
rect 68348 81678 68350 81730
rect 68402 81678 68404 81730
rect 68348 81284 68404 81678
rect 68460 81284 68516 81294
rect 68348 81282 68516 81284
rect 68348 81230 68462 81282
rect 68514 81230 68516 81282
rect 68348 81228 68516 81230
rect 68460 81218 68516 81228
rect 68572 80498 68628 80510
rect 68572 80446 68574 80498
rect 68626 80446 68628 80498
rect 68572 80276 68628 80446
rect 68572 80210 68628 80220
rect 68236 80098 68292 80108
rect 68124 79550 68126 79602
rect 68178 79550 68180 79602
rect 68124 78988 68180 79550
rect 68684 79602 68740 82236
rect 69244 82292 69300 84142
rect 69356 83410 69412 88844
rect 70476 88002 70532 88844
rect 71036 88898 71092 88910
rect 71036 88846 71038 88898
rect 71090 88846 71092 88898
rect 71036 88228 71092 88846
rect 71596 88900 71652 88910
rect 71596 88806 71652 88844
rect 70476 87950 70478 88002
rect 70530 87950 70532 88002
rect 70252 87330 70308 87342
rect 70252 87278 70254 87330
rect 70306 87278 70308 87330
rect 69804 86660 69860 86670
rect 69804 86566 69860 86604
rect 70252 86660 70308 87278
rect 70252 86594 70308 86604
rect 70140 86546 70196 86558
rect 70140 86494 70142 86546
rect 70194 86494 70196 86546
rect 69468 86436 69524 86446
rect 69468 86342 69524 86380
rect 70140 86324 70196 86494
rect 70364 86546 70420 86558
rect 70364 86494 70366 86546
rect 70418 86494 70420 86546
rect 70364 86436 70420 86494
rect 70364 86370 70420 86380
rect 70140 86258 70196 86268
rect 70364 86100 70420 86110
rect 69356 83358 69358 83410
rect 69410 83358 69412 83410
rect 69356 83346 69412 83358
rect 69468 85764 69524 85774
rect 69468 85090 69524 85708
rect 69468 85038 69470 85090
rect 69522 85038 69524 85090
rect 69244 82226 69300 82236
rect 69468 82626 69524 85038
rect 70140 84980 70196 84990
rect 70140 84978 70308 84980
rect 70140 84926 70142 84978
rect 70194 84926 70308 84978
rect 70140 84924 70308 84926
rect 70140 84914 70196 84924
rect 70140 84084 70196 84094
rect 69692 84082 70196 84084
rect 69692 84030 70142 84082
rect 70194 84030 70196 84082
rect 69692 84028 70196 84030
rect 69692 83522 69748 84028
rect 70140 84018 70196 84028
rect 69692 83470 69694 83522
rect 69746 83470 69748 83522
rect 69692 83458 69748 83470
rect 70252 83410 70308 84924
rect 70364 84084 70420 86044
rect 70476 85764 70532 87950
rect 70588 88172 71092 88228
rect 70588 86436 70644 88172
rect 71036 88002 71092 88014
rect 71036 87950 71038 88002
rect 71090 87950 71092 88002
rect 71036 87556 71092 87950
rect 71932 87892 71988 87902
rect 71036 87500 71540 87556
rect 70588 86370 70644 86380
rect 70700 87442 70756 87454
rect 70700 87390 70702 87442
rect 70754 87390 70756 87442
rect 70700 86324 70756 87390
rect 71372 87220 71428 87230
rect 70700 86258 70756 86268
rect 70812 87218 71428 87220
rect 70812 87166 71374 87218
rect 71426 87166 71428 87218
rect 70812 87164 71428 87166
rect 71484 87220 71540 87500
rect 71932 87444 71988 87836
rect 71708 87220 71764 87230
rect 71484 87218 71764 87220
rect 71484 87166 71710 87218
rect 71762 87166 71764 87218
rect 71484 87164 71764 87166
rect 70476 85698 70532 85708
rect 70812 85316 70868 87164
rect 71372 87154 71428 87164
rect 71372 86548 71428 86558
rect 71372 86454 71428 86492
rect 70588 85260 70868 85316
rect 71036 86436 71092 86446
rect 70476 84084 70532 84094
rect 70364 84082 70532 84084
rect 70364 84030 70478 84082
rect 70530 84030 70532 84082
rect 70364 84028 70532 84030
rect 70252 83358 70254 83410
rect 70306 83358 70308 83410
rect 70252 83346 70308 83358
rect 69468 82574 69470 82626
rect 69522 82574 69524 82626
rect 69468 81396 69524 82574
rect 69916 82628 69972 82638
rect 70476 82628 70532 84028
rect 70588 83522 70644 85260
rect 71036 84418 71092 86380
rect 71596 86100 71652 87164
rect 71708 87154 71764 87164
rect 71596 86034 71652 86044
rect 71708 86660 71764 86670
rect 71036 84366 71038 84418
rect 71090 84366 71092 84418
rect 71036 84354 71092 84366
rect 71708 85762 71764 86604
rect 71932 86546 71988 87388
rect 71932 86494 71934 86546
rect 71986 86494 71988 86546
rect 71932 86482 71988 86494
rect 72268 87554 72324 87566
rect 72268 87502 72270 87554
rect 72322 87502 72324 87554
rect 72268 86546 72324 87502
rect 72492 87442 72548 87454
rect 72492 87390 72494 87442
rect 72546 87390 72548 87442
rect 72492 87332 72548 87390
rect 72492 87266 72548 87276
rect 73164 87444 73220 87454
rect 73164 87332 73220 87388
rect 73276 87332 73332 87342
rect 73164 87330 73332 87332
rect 73164 87278 73278 87330
rect 73330 87278 73332 87330
rect 73164 87276 73332 87278
rect 73164 86770 73220 87276
rect 73276 87266 73332 87276
rect 73724 87332 73780 87342
rect 74508 87332 74564 87342
rect 75068 87332 75124 87342
rect 75516 87332 75572 87342
rect 73780 87276 73892 87332
rect 73724 87200 73780 87276
rect 73164 86718 73166 86770
rect 73218 86718 73220 86770
rect 73164 86706 73220 86718
rect 72268 86494 72270 86546
rect 72322 86494 72324 86546
rect 71708 85710 71710 85762
rect 71762 85710 71764 85762
rect 70588 83470 70590 83522
rect 70642 83470 70644 83522
rect 70588 83458 70644 83470
rect 71260 84306 71316 84318
rect 71260 84254 71262 84306
rect 71314 84254 71316 84306
rect 71260 83300 71316 84254
rect 71260 83234 71316 83244
rect 71596 83300 71652 83310
rect 71596 83206 71652 83244
rect 69916 82626 70532 82628
rect 69916 82574 69918 82626
rect 69970 82574 70532 82626
rect 69916 82572 70532 82574
rect 69804 81732 69860 81742
rect 69468 81330 69524 81340
rect 69580 81730 69860 81732
rect 69580 81678 69806 81730
rect 69858 81678 69860 81730
rect 69580 81676 69860 81678
rect 69244 81170 69300 81182
rect 69244 81118 69246 81170
rect 69298 81118 69300 81170
rect 69244 80612 69300 81118
rect 69244 80546 69300 80556
rect 69468 80276 69524 80286
rect 69468 80182 69524 80220
rect 69580 80274 69636 81676
rect 69804 81666 69860 81676
rect 69692 81396 69748 81406
rect 69692 81302 69748 81340
rect 69580 80222 69582 80274
rect 69634 80222 69636 80274
rect 69244 80164 69300 80174
rect 69244 80070 69300 80108
rect 69580 80052 69636 80222
rect 69580 79828 69636 79996
rect 69580 79762 69636 79772
rect 69692 80948 69748 80958
rect 68684 79550 68686 79602
rect 68738 79550 68740 79602
rect 68684 79538 68740 79550
rect 69580 79604 69636 79614
rect 69692 79604 69748 80892
rect 69580 79602 69748 79604
rect 69580 79550 69582 79602
rect 69634 79550 69748 79602
rect 69580 79548 69748 79550
rect 69580 79538 69636 79548
rect 67676 78932 68180 78988
rect 67676 78372 67732 78932
rect 68572 78820 68628 78830
rect 67900 78818 68628 78820
rect 67900 78766 68574 78818
rect 68626 78766 68628 78818
rect 67900 78764 68628 78766
rect 67676 78258 67732 78316
rect 67676 78206 67678 78258
rect 67730 78206 67732 78258
rect 67676 78194 67732 78206
rect 67788 78708 67844 78718
rect 67788 78260 67844 78652
rect 67788 78194 67844 78204
rect 67900 78706 67956 78764
rect 68572 78754 68628 78764
rect 69580 78818 69636 78830
rect 69580 78766 69582 78818
rect 69634 78766 69636 78818
rect 67900 78654 67902 78706
rect 67954 78654 67956 78706
rect 67900 77476 67956 78654
rect 69020 78708 69076 78718
rect 68124 78594 68180 78606
rect 68124 78542 68126 78594
rect 68178 78542 68180 78594
rect 68124 78260 68180 78542
rect 68124 78194 68180 78204
rect 69020 78146 69076 78652
rect 69020 78094 69022 78146
rect 69074 78094 69076 78146
rect 68012 78036 68068 78046
rect 68460 78036 68516 78046
rect 68012 78034 68516 78036
rect 68012 77982 68014 78034
rect 68066 77982 68462 78034
rect 68514 77982 68516 78034
rect 68012 77980 68516 77982
rect 68012 77970 68068 77980
rect 67788 77420 67956 77476
rect 68460 77476 68516 77980
rect 67788 76692 67844 77420
rect 67900 77252 67956 77262
rect 67900 77158 67956 77196
rect 68348 77028 68404 77038
rect 67788 76020 67844 76636
rect 68236 77026 68404 77028
rect 68236 76974 68350 77026
rect 68402 76974 68404 77026
rect 68236 76972 68404 76974
rect 68124 76468 68180 76478
rect 68124 76374 68180 76412
rect 67788 75954 67844 75964
rect 67564 75906 67620 75918
rect 67564 75854 67566 75906
rect 67618 75854 67620 75906
rect 67564 75794 67620 75854
rect 68124 75908 68180 75918
rect 68236 75908 68292 76972
rect 68348 76962 68404 76972
rect 68460 76804 68516 77420
rect 69020 77364 69076 78094
rect 69356 78596 69412 78606
rect 69356 78146 69412 78540
rect 69356 78094 69358 78146
rect 69410 78094 69412 78146
rect 69356 78082 69412 78094
rect 69244 77364 69300 77374
rect 69020 77362 69300 77364
rect 69020 77310 69246 77362
rect 69298 77310 69300 77362
rect 69020 77308 69300 77310
rect 69244 77298 69300 77308
rect 68124 75906 68292 75908
rect 68124 75854 68126 75906
rect 68178 75854 68292 75906
rect 68124 75852 68292 75854
rect 68348 76748 68516 76804
rect 69580 77252 69636 78766
rect 69804 78820 69860 78830
rect 69804 78258 69860 78764
rect 69804 78206 69806 78258
rect 69858 78206 69860 78258
rect 69804 78194 69860 78206
rect 69580 77028 69636 77196
rect 69692 77028 69748 77038
rect 69580 77026 69748 77028
rect 69580 76974 69694 77026
rect 69746 76974 69748 77026
rect 69580 76972 69748 76974
rect 68124 75842 68180 75852
rect 67564 75742 67566 75794
rect 67618 75742 67620 75794
rect 67564 74226 67620 75742
rect 68012 75684 68068 75694
rect 68012 75590 68068 75628
rect 67788 74788 67844 74798
rect 67788 74786 68292 74788
rect 67788 74734 67790 74786
rect 67842 74734 68292 74786
rect 67788 74732 68292 74734
rect 67788 74722 67844 74732
rect 67564 74174 67566 74226
rect 67618 74174 67620 74226
rect 67564 73556 67620 74174
rect 67564 73490 67620 73500
rect 68236 73554 68292 74732
rect 68236 73502 68238 73554
rect 68290 73502 68292 73554
rect 68236 73490 68292 73502
rect 68012 71652 68068 71662
rect 68012 71650 68292 71652
rect 68012 71598 68014 71650
rect 68066 71598 68292 71650
rect 68012 71596 68292 71598
rect 68012 71586 68068 71596
rect 68124 71092 68180 71102
rect 67452 70466 67508 70476
rect 67788 70754 67844 70766
rect 67788 70702 67790 70754
rect 67842 70702 67844 70754
rect 67788 70308 67844 70702
rect 67340 70306 67732 70308
rect 67340 70254 67342 70306
rect 67394 70254 67732 70306
rect 67340 70252 67732 70254
rect 67340 70242 67396 70252
rect 66556 69970 66612 69982
rect 66556 69918 66558 69970
rect 66610 69918 66612 69970
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 65548 68850 66164 68852
rect 65548 68798 65550 68850
rect 65602 68798 66164 68850
rect 65548 68796 66164 68798
rect 65548 68786 65604 68796
rect 66108 68626 66164 68796
rect 66108 68574 66110 68626
rect 66162 68574 66164 68626
rect 66108 68562 66164 68574
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 66556 67620 66612 69918
rect 67676 69524 67732 70252
rect 67788 70242 67844 70252
rect 68124 70194 68180 71036
rect 68236 70866 68292 71596
rect 68236 70814 68238 70866
rect 68290 70814 68292 70866
rect 68236 70756 68292 70814
rect 68236 70690 68292 70700
rect 68124 70142 68126 70194
rect 68178 70142 68180 70194
rect 68124 70130 68180 70142
rect 67564 69298 67620 69310
rect 67564 69246 67566 69298
rect 67618 69246 67620 69298
rect 67340 69188 67396 69198
rect 66892 68514 66948 68526
rect 66892 68462 66894 68514
rect 66946 68462 66948 68514
rect 66892 67844 66948 68462
rect 67228 68292 67284 68302
rect 66892 67778 66948 67788
rect 67004 67954 67060 67966
rect 67004 67902 67006 67954
rect 67058 67902 67060 67954
rect 67004 67620 67060 67902
rect 66332 67564 67060 67620
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65996 66500 66052 66510
rect 66332 66500 66388 67564
rect 66556 67060 66612 67070
rect 65996 66498 66388 66500
rect 65996 66446 65998 66498
rect 66050 66446 66388 66498
rect 65996 66444 66388 66446
rect 66444 67058 66612 67060
rect 66444 67006 66558 67058
rect 66610 67006 66612 67058
rect 66444 67004 66612 67006
rect 65996 66434 66052 66444
rect 65436 65650 65492 65660
rect 65660 66050 65716 66062
rect 65660 65998 65662 66050
rect 65714 65998 65716 66050
rect 65660 65604 65716 65998
rect 65660 65538 65716 65548
rect 66332 65604 66388 65614
rect 66444 65604 66500 67004
rect 66556 66994 66612 67004
rect 66332 65602 66500 65604
rect 66332 65550 66334 65602
rect 66386 65550 66500 65602
rect 66332 65548 66500 65550
rect 66556 66276 66612 66286
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 66332 64708 66388 65548
rect 66556 64820 66612 66220
rect 66780 66162 66836 66174
rect 66780 66110 66782 66162
rect 66834 66110 66836 66162
rect 66220 64148 66276 64158
rect 66220 64054 66276 64092
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 66220 63364 66276 63374
rect 66220 63250 66276 63308
rect 66220 63198 66222 63250
rect 66274 63198 66276 63250
rect 66220 63186 66276 63198
rect 65884 62916 65940 62926
rect 65884 62822 65940 62860
rect 66332 62354 66388 64652
rect 66332 62302 66334 62354
rect 66386 62302 66388 62354
rect 66332 62290 66388 62302
rect 66444 64764 66612 64820
rect 66668 65492 66724 65502
rect 65772 62244 65828 62282
rect 65324 62132 65492 62188
rect 65772 62178 65828 62188
rect 64876 60564 64932 60574
rect 64876 59890 64932 60508
rect 64876 59838 64878 59890
rect 64930 59838 64932 59890
rect 64876 59826 64932 59838
rect 65100 60002 65156 62132
rect 65324 60900 65380 60910
rect 65324 60806 65380 60844
rect 65100 59950 65102 60002
rect 65154 59950 65156 60002
rect 65100 59892 65156 59950
rect 65100 59826 65156 59836
rect 64428 59724 64820 59780
rect 64204 58436 64260 58446
rect 64204 58342 64260 58380
rect 64316 58212 64372 58222
rect 64316 56978 64372 58156
rect 64316 56926 64318 56978
rect 64370 56926 64372 56978
rect 64316 56914 64372 56926
rect 64316 54740 64372 54750
rect 64204 54628 64260 54638
rect 64204 54534 64260 54572
rect 64316 54626 64372 54684
rect 64316 54574 64318 54626
rect 64370 54574 64372 54626
rect 64316 54562 64372 54574
rect 64316 53842 64372 53854
rect 64316 53790 64318 53842
rect 64370 53790 64372 53842
rect 64316 53172 64372 53790
rect 64316 53106 64372 53116
rect 63980 51602 64092 51604
rect 63980 51550 63982 51602
rect 64034 51550 64092 51602
rect 63980 51548 64092 51550
rect 63980 51538 64036 51548
rect 64092 51538 64148 51548
rect 64092 51380 64148 51390
rect 64092 51286 64148 51324
rect 63980 51156 64036 51166
rect 63868 51154 64036 51156
rect 63868 51102 63982 51154
rect 64034 51102 64036 51154
rect 63868 51100 64036 51102
rect 63868 50428 63924 51100
rect 63980 51090 64036 51100
rect 63532 50372 63924 50428
rect 63420 48354 63476 48366
rect 63420 48302 63422 48354
rect 63474 48302 63476 48354
rect 63420 48132 63476 48302
rect 63532 48354 63588 50372
rect 64204 48468 64260 48478
rect 64204 48374 64260 48412
rect 63532 48302 63534 48354
rect 63586 48302 63588 48354
rect 63532 48290 63588 48302
rect 64316 48244 64372 48254
rect 64316 48150 64372 48188
rect 63420 48066 63476 48076
rect 64204 48020 64260 48030
rect 64204 47926 64260 47964
rect 64204 47124 64260 47134
rect 64204 46004 64260 47068
rect 64316 46788 64372 46798
rect 64316 46562 64372 46732
rect 64316 46510 64318 46562
rect 64370 46510 64372 46562
rect 64316 46498 64372 46510
rect 64316 46004 64372 46014
rect 64204 46002 64372 46004
rect 64204 45950 64318 46002
rect 64370 45950 64372 46002
rect 64204 45948 64372 45950
rect 64316 45938 64372 45948
rect 63532 45444 63588 45454
rect 63532 45218 63588 45388
rect 63532 45166 63534 45218
rect 63586 45166 63588 45218
rect 63532 45154 63588 45166
rect 64204 45106 64260 45118
rect 64204 45054 64206 45106
rect 64258 45054 64260 45106
rect 63420 43764 63476 43774
rect 63420 43670 63476 43708
rect 64204 43652 64260 45054
rect 64428 44548 64484 59724
rect 65436 59556 65492 62132
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65996 61684 66052 61694
rect 65996 61590 66052 61628
rect 65548 61346 65604 61358
rect 65548 61294 65550 61346
rect 65602 61294 65604 61346
rect 65548 60900 65604 61294
rect 65548 60834 65604 60844
rect 66220 61124 66276 61134
rect 65884 60788 65940 60798
rect 65884 60674 65940 60732
rect 65884 60622 65886 60674
rect 65938 60622 65940 60674
rect 65884 60562 65940 60622
rect 66220 60676 66276 61068
rect 66444 60788 66500 64764
rect 66668 64034 66724 65436
rect 66668 63982 66670 64034
rect 66722 63982 66724 64034
rect 66668 63924 66724 63982
rect 66668 63858 66724 63868
rect 66780 64820 66836 66110
rect 67004 65828 67060 65838
rect 66892 64820 66948 64830
rect 66780 64818 66948 64820
rect 66780 64766 66894 64818
rect 66946 64766 66948 64818
rect 66780 64764 66948 64766
rect 66556 63364 66612 63374
rect 66556 61684 66612 63308
rect 66556 61570 66612 61628
rect 66556 61518 66558 61570
rect 66610 61518 66612 61570
rect 66556 61506 66612 61518
rect 66668 61012 66724 61022
rect 66668 60918 66724 60956
rect 66444 60732 66724 60788
rect 66220 60674 66388 60676
rect 66220 60622 66222 60674
rect 66274 60622 66388 60674
rect 66220 60620 66388 60622
rect 66220 60610 66276 60620
rect 65884 60510 65886 60562
rect 65938 60510 65940 60562
rect 65884 60498 65940 60510
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 66108 60226 66164 60238
rect 66108 60174 66110 60226
rect 66162 60174 66164 60226
rect 65548 60002 65604 60014
rect 65548 59950 65550 60002
rect 65602 59950 65604 60002
rect 65548 59780 65604 59950
rect 65884 59892 65940 59902
rect 65548 59714 65604 59724
rect 65660 59890 65940 59892
rect 65660 59838 65886 59890
rect 65938 59838 65940 59890
rect 65660 59836 65940 59838
rect 65436 59490 65492 59500
rect 65324 59220 65380 59230
rect 64540 59106 64596 59118
rect 64540 59054 64542 59106
rect 64594 59054 64596 59106
rect 64540 58436 64596 59054
rect 64988 58660 65044 58670
rect 64988 58566 65044 58604
rect 65100 58436 65156 58446
rect 64596 58380 64708 58436
rect 64540 58370 64596 58380
rect 64540 55970 64596 55982
rect 64540 55918 64542 55970
rect 64594 55918 64596 55970
rect 64540 53844 64596 55918
rect 64540 53778 64596 53788
rect 64652 53732 64708 58380
rect 65100 58342 65156 58380
rect 64988 58212 65044 58222
rect 64988 58118 65044 58156
rect 65324 57874 65380 59164
rect 65548 58324 65604 58334
rect 65548 58230 65604 58268
rect 65660 58212 65716 59836
rect 65884 59826 65940 59836
rect 65884 59220 65940 59230
rect 66108 59220 66164 60174
rect 66332 60228 66388 60620
rect 66556 60562 66612 60574
rect 66556 60510 66558 60562
rect 66610 60510 66612 60562
rect 66332 60172 66500 60228
rect 66332 59780 66388 59790
rect 66332 59686 66388 59724
rect 65884 59218 66164 59220
rect 65884 59166 65886 59218
rect 65938 59166 66164 59218
rect 65884 59164 66164 59166
rect 66444 59220 66500 60172
rect 66556 59332 66612 60510
rect 66668 59668 66724 60732
rect 66780 60226 66836 64764
rect 66892 64754 66948 64764
rect 67004 64036 67060 65772
rect 67004 63922 67060 63980
rect 67004 63870 67006 63922
rect 67058 63870 67060 63922
rect 67004 63858 67060 63870
rect 66892 62916 66948 62926
rect 66892 61346 66948 62860
rect 67116 62916 67172 62926
rect 67116 62822 67172 62860
rect 66892 61294 66894 61346
rect 66946 61294 66948 61346
rect 66892 60564 66948 61294
rect 67116 62242 67172 62254
rect 67116 62190 67118 62242
rect 67170 62190 67172 62242
rect 67116 60788 67172 62190
rect 67228 61348 67284 68236
rect 67340 67170 67396 69132
rect 67564 68516 67620 69246
rect 67676 69298 67732 69468
rect 67676 69246 67678 69298
rect 67730 69246 67732 69298
rect 67676 69234 67732 69246
rect 67900 69188 67956 69198
rect 67452 67844 67508 67854
rect 67452 67750 67508 67788
rect 67564 67620 67620 68460
rect 67788 69186 67956 69188
rect 67788 69134 67902 69186
rect 67954 69134 67956 69186
rect 67788 69132 67956 69134
rect 67788 68068 67844 69132
rect 67900 69122 67956 69132
rect 68236 69188 68292 69198
rect 68236 69094 68292 69132
rect 68348 68292 68404 76748
rect 68908 76356 68964 76366
rect 68908 76354 69412 76356
rect 68908 76302 68910 76354
rect 68962 76302 69412 76354
rect 68908 76300 69412 76302
rect 68908 76290 68964 76300
rect 69356 75570 69412 76300
rect 69356 75518 69358 75570
rect 69410 75518 69412 75570
rect 69356 75506 69412 75518
rect 68572 74004 68628 74014
rect 68572 73442 68628 73948
rect 69468 74004 69524 74014
rect 69468 73910 69524 73948
rect 68572 73390 68574 73442
rect 68626 73390 68628 73442
rect 68572 73378 68628 73390
rect 69244 72324 69300 72334
rect 69580 72324 69636 76972
rect 69692 76962 69748 76972
rect 69916 75796 69972 82572
rect 70364 81732 70420 81742
rect 70364 81730 70532 81732
rect 70364 81678 70366 81730
rect 70418 81678 70532 81730
rect 70364 81676 70532 81678
rect 70364 81666 70420 81676
rect 70140 81060 70196 81070
rect 70140 80966 70196 81004
rect 70476 80612 70532 81676
rect 71484 81172 71540 81182
rect 71372 81116 71484 81172
rect 70588 81058 70644 81070
rect 70588 81006 70590 81058
rect 70642 81006 70644 81058
rect 70588 80948 70644 81006
rect 70588 80882 70644 80892
rect 71148 81058 71204 81070
rect 71148 81006 71150 81058
rect 71202 81006 71204 81058
rect 71148 80946 71204 81006
rect 71148 80894 71150 80946
rect 71202 80894 71204 80946
rect 71148 80882 71204 80894
rect 70028 80388 70084 80398
rect 70028 80294 70084 80332
rect 70364 80388 70420 80398
rect 70364 80294 70420 80332
rect 70140 80164 70196 80174
rect 70028 78260 70084 78270
rect 70028 78166 70084 78204
rect 70140 78146 70196 80108
rect 70252 80162 70308 80174
rect 70252 80110 70254 80162
rect 70306 80110 70308 80162
rect 70252 79716 70308 80110
rect 70252 79650 70308 79660
rect 70364 80164 70420 80174
rect 70476 80164 70532 80556
rect 70420 80108 70532 80164
rect 70700 80500 70756 80510
rect 70364 78988 70420 80108
rect 70700 79828 70756 80444
rect 71372 80388 71428 81116
rect 71484 81078 71540 81116
rect 70812 80276 70868 80286
rect 70812 80182 70868 80220
rect 70812 79828 70868 79838
rect 70700 79826 70868 79828
rect 70700 79774 70814 79826
rect 70866 79774 70868 79826
rect 70700 79772 70868 79774
rect 70476 79604 70532 79614
rect 70476 79602 70756 79604
rect 70476 79550 70478 79602
rect 70530 79550 70756 79602
rect 70476 79548 70756 79550
rect 70476 79538 70532 79548
rect 70700 78988 70756 79548
rect 70364 78932 70532 78988
rect 70140 78094 70142 78146
rect 70194 78094 70196 78146
rect 70140 78082 70196 78094
rect 70476 78036 70532 78932
rect 70588 78932 70756 78988
rect 70588 78596 70644 78932
rect 70588 78258 70644 78540
rect 70588 78206 70590 78258
rect 70642 78206 70644 78258
rect 70588 78194 70644 78206
rect 70476 77980 70644 78036
rect 70588 76468 70644 77980
rect 70812 77252 70868 79772
rect 71372 79826 71428 80332
rect 71596 80946 71652 80958
rect 71596 80894 71598 80946
rect 71650 80894 71652 80946
rect 71372 79774 71374 79826
rect 71426 79774 71428 79826
rect 71372 79762 71428 79774
rect 71484 80276 71540 80286
rect 71484 79604 71540 80220
rect 71484 78036 71540 79548
rect 71596 79602 71652 80894
rect 71708 80948 71764 85710
rect 71932 86324 71988 86334
rect 71932 84306 71988 86268
rect 72268 85202 72324 86494
rect 73388 86660 73444 86670
rect 72716 86100 72772 86110
rect 72716 86006 72772 86044
rect 73388 86100 73444 86604
rect 73724 86660 73780 86670
rect 73724 86566 73780 86604
rect 73388 85968 73444 86044
rect 73836 85764 73892 87276
rect 74508 87330 74788 87332
rect 74508 87278 74510 87330
rect 74562 87278 74788 87330
rect 74508 87276 74788 87278
rect 74508 87266 74564 87276
rect 74732 86772 74788 87276
rect 75068 87330 75572 87332
rect 75068 87278 75070 87330
rect 75122 87278 75518 87330
rect 75570 87278 75572 87330
rect 75068 87276 75572 87278
rect 75068 87266 75124 87276
rect 74732 86770 74900 86772
rect 74732 86718 74734 86770
rect 74786 86718 74900 86770
rect 74732 86716 74900 86718
rect 74732 86706 74788 86716
rect 74396 86660 74452 86670
rect 74396 86566 74452 86604
rect 74620 85874 74676 85886
rect 74620 85822 74622 85874
rect 74674 85822 74676 85874
rect 73836 85762 74004 85764
rect 73836 85710 73838 85762
rect 73890 85710 74004 85762
rect 73836 85708 74004 85710
rect 73836 85698 73892 85708
rect 72268 85150 72270 85202
rect 72322 85150 72324 85202
rect 72268 85138 72324 85150
rect 73164 85652 73220 85662
rect 73164 85202 73220 85596
rect 73164 85150 73166 85202
rect 73218 85150 73220 85202
rect 73164 85138 73220 85150
rect 72828 84866 72884 84878
rect 72828 84814 72830 84866
rect 72882 84814 72884 84866
rect 71932 84254 71934 84306
rect 71986 84254 71988 84306
rect 71932 84242 71988 84254
rect 72492 84308 72548 84318
rect 72828 84308 72884 84814
rect 73948 84532 74004 85708
rect 74060 85092 74116 85102
rect 74060 85090 74228 85092
rect 74060 85038 74062 85090
rect 74114 85038 74228 85090
rect 74060 85036 74228 85038
rect 74060 85026 74116 85036
rect 73948 84466 74004 84476
rect 72492 84306 72884 84308
rect 72492 84254 72494 84306
rect 72546 84254 72884 84306
rect 72492 84252 72884 84254
rect 73612 84308 73668 84318
rect 72492 83524 72548 84252
rect 73612 84214 73668 84252
rect 74172 83748 74228 85036
rect 74284 84866 74340 84878
rect 74284 84814 74286 84866
rect 74338 84814 74340 84866
rect 74284 84418 74340 84814
rect 74284 84366 74286 84418
rect 74338 84366 74340 84418
rect 74284 84354 74340 84366
rect 74620 84308 74676 85822
rect 74620 84242 74676 84252
rect 74732 85764 74788 85774
rect 74284 83748 74340 83758
rect 74172 83746 74340 83748
rect 74172 83694 74286 83746
rect 74338 83694 74340 83746
rect 74172 83692 74340 83694
rect 74284 83682 74340 83692
rect 74620 83748 74676 83758
rect 74732 83748 74788 85708
rect 74844 84980 74900 86716
rect 75516 86660 75572 87276
rect 74956 86548 75012 86558
rect 74956 85314 75012 86492
rect 75404 86434 75460 86446
rect 75404 86382 75406 86434
rect 75458 86382 75460 86434
rect 75292 85988 75348 85998
rect 75404 85988 75460 86382
rect 75292 85986 75460 85988
rect 75292 85934 75294 85986
rect 75346 85934 75460 85986
rect 75292 85932 75460 85934
rect 75292 85922 75348 85932
rect 74956 85262 74958 85314
rect 75010 85262 75012 85314
rect 74956 85250 75012 85262
rect 75292 85764 75348 85774
rect 75516 85764 75572 86604
rect 77868 86658 77924 86670
rect 77868 86606 77870 86658
rect 77922 86606 77924 86658
rect 75740 86548 75796 86558
rect 75740 86454 75796 86492
rect 76524 86434 76580 86446
rect 76524 86382 76526 86434
rect 76578 86382 76580 86434
rect 76524 85876 76580 86382
rect 76524 85810 76580 85820
rect 77308 86434 77364 86446
rect 77308 86382 77310 86434
rect 77362 86382 77364 86434
rect 76076 85764 76132 85774
rect 75516 85708 75796 85764
rect 75292 85314 75348 85708
rect 75292 85262 75294 85314
rect 75346 85262 75348 85314
rect 75292 85250 75348 85262
rect 74844 84914 74900 84924
rect 75628 84980 75684 84990
rect 75628 84886 75684 84924
rect 75516 84308 75572 84318
rect 74620 83746 74788 83748
rect 74620 83694 74622 83746
rect 74674 83694 74788 83746
rect 74620 83692 74788 83694
rect 74620 83682 74676 83692
rect 72716 83524 72772 83534
rect 72492 83522 72772 83524
rect 72492 83470 72718 83522
rect 72770 83470 72772 83522
rect 72492 83468 72772 83470
rect 72716 81844 72772 83468
rect 73164 83522 73220 83534
rect 73164 83470 73166 83522
rect 73218 83470 73220 83522
rect 73164 83300 73220 83470
rect 73164 83234 73220 83244
rect 73612 83298 73668 83310
rect 73612 83246 73614 83298
rect 73666 83246 73668 83298
rect 73276 82628 73332 82638
rect 73276 82066 73332 82572
rect 73276 82014 73278 82066
rect 73330 82014 73332 82066
rect 72828 81844 72884 81854
rect 72716 81788 72828 81844
rect 72828 81750 72884 81788
rect 73276 81732 73332 82014
rect 73612 81844 73668 83246
rect 74732 82964 74788 83692
rect 75404 84084 75460 84094
rect 74956 83410 75012 83422
rect 74956 83358 74958 83410
rect 75010 83358 75012 83410
rect 74844 82964 74900 82974
rect 74732 82962 74900 82964
rect 74732 82910 74846 82962
rect 74898 82910 74900 82962
rect 74732 82908 74900 82910
rect 73836 82628 73892 82638
rect 73836 82534 73892 82572
rect 74844 81956 74900 82908
rect 74956 82628 75012 83358
rect 75404 83410 75460 84028
rect 75404 83358 75406 83410
rect 75458 83358 75460 83410
rect 75404 83346 75460 83358
rect 75516 82738 75572 84252
rect 75516 82686 75518 82738
rect 75570 82686 75572 82738
rect 75516 82674 75572 82686
rect 74956 82562 75012 82572
rect 75404 82068 75460 82078
rect 75404 81974 75460 82012
rect 74844 81900 75236 81956
rect 73612 81778 73668 81788
rect 73276 81666 73332 81676
rect 73836 81732 73892 81742
rect 73836 81638 73892 81676
rect 74284 81732 74340 81742
rect 74284 81638 74340 81676
rect 74844 81732 74900 81742
rect 73836 81396 73892 81406
rect 73836 81302 73892 81340
rect 74508 81396 74564 81406
rect 74508 81394 74788 81396
rect 74508 81342 74510 81394
rect 74562 81342 74788 81394
rect 74508 81340 74788 81342
rect 74508 81330 74564 81340
rect 72604 81172 72660 81182
rect 73500 81172 73556 81182
rect 72268 81170 73556 81172
rect 72268 81118 72606 81170
rect 72658 81118 73502 81170
rect 73554 81118 73556 81170
rect 72268 81116 73556 81118
rect 71708 80882 71764 80892
rect 72044 81058 72100 81070
rect 72044 81006 72046 81058
rect 72098 81006 72100 81058
rect 72044 80946 72100 81006
rect 72044 80894 72046 80946
rect 72098 80894 72100 80946
rect 72044 80882 72100 80894
rect 71708 80386 71764 80398
rect 71708 80334 71710 80386
rect 71762 80334 71764 80386
rect 71708 80164 71764 80334
rect 71708 80098 71764 80108
rect 72268 80052 72324 81116
rect 72604 81106 72660 81116
rect 73500 81106 73556 81116
rect 74284 81170 74340 81182
rect 74284 81118 74286 81170
rect 74338 81118 74340 81170
rect 72380 80276 72436 80286
rect 72380 80274 72884 80276
rect 72380 80222 72382 80274
rect 72434 80222 72884 80274
rect 72380 80220 72884 80222
rect 72380 80210 72436 80220
rect 72268 79996 72548 80052
rect 72268 79828 72324 79838
rect 72268 79734 72324 79772
rect 71596 79550 71598 79602
rect 71650 79550 71652 79602
rect 71596 78988 71652 79550
rect 72492 79602 72548 79996
rect 72492 79550 72494 79602
rect 72546 79550 72548 79602
rect 72492 78988 72548 79550
rect 71596 78932 71764 78988
rect 72492 78932 72660 78988
rect 71708 78708 71764 78932
rect 71708 78642 71764 78652
rect 71596 78036 71652 78046
rect 71484 78034 71652 78036
rect 71484 77982 71598 78034
rect 71650 77982 71652 78034
rect 71484 77980 71652 77982
rect 71596 77970 71652 77980
rect 72044 78034 72100 78046
rect 72044 77982 72046 78034
rect 72098 77982 72100 78034
rect 71036 77924 71092 77934
rect 71036 77922 71204 77924
rect 71036 77870 71038 77922
rect 71090 77870 71204 77922
rect 71036 77868 71204 77870
rect 71036 77858 71092 77868
rect 70812 77120 70868 77196
rect 70140 75796 70196 75806
rect 69916 75794 70532 75796
rect 69916 75742 70142 75794
rect 70194 75742 70532 75794
rect 69916 75740 70532 75742
rect 70140 75730 70196 75740
rect 69692 75570 69748 75582
rect 69692 75518 69694 75570
rect 69746 75518 69748 75570
rect 69692 75124 69748 75518
rect 70476 75348 70532 75740
rect 70588 75794 70644 76412
rect 70588 75742 70590 75794
rect 70642 75742 70644 75794
rect 70588 75730 70644 75742
rect 71036 76354 71092 76366
rect 71036 76302 71038 76354
rect 71090 76302 71092 76354
rect 70476 75292 70980 75348
rect 69692 75058 69748 75068
rect 70588 75124 70644 75134
rect 70588 75030 70644 75068
rect 70924 74900 70980 75292
rect 71036 75012 71092 76302
rect 71148 75796 71204 77868
rect 71820 77252 71876 77262
rect 71820 77158 71876 77196
rect 71260 77026 71316 77038
rect 71260 76974 71262 77026
rect 71314 76974 71316 77026
rect 71260 76468 71316 76974
rect 71932 77026 71988 77038
rect 71932 76974 71934 77026
rect 71986 76974 71988 77026
rect 71260 76402 71316 76412
rect 71596 76466 71652 76478
rect 71596 76414 71598 76466
rect 71650 76414 71652 76466
rect 71260 75796 71316 75806
rect 71148 75740 71260 75796
rect 71260 75702 71316 75740
rect 71596 75796 71652 76414
rect 71932 76356 71988 76974
rect 71932 76290 71988 76300
rect 71596 75730 71652 75740
rect 72044 75796 72100 77982
rect 72604 77924 72660 78932
rect 72604 77858 72660 77868
rect 72828 77474 72884 80220
rect 73836 80164 73892 80174
rect 73500 79602 73556 79614
rect 73500 79550 73502 79602
rect 73554 79550 73556 79602
rect 73500 78036 73556 79550
rect 73836 78930 73892 80108
rect 74172 79716 74228 79726
rect 74284 79716 74340 81118
rect 74620 81170 74676 81182
rect 74620 81118 74622 81170
rect 74674 81118 74676 81170
rect 74620 80724 74676 81118
rect 74396 80668 74676 80724
rect 74732 80724 74788 81340
rect 74844 81172 74900 81676
rect 75180 81620 75236 81900
rect 75740 81732 75796 85708
rect 76076 84978 76132 85708
rect 76076 84926 76078 84978
rect 76130 84926 76132 84978
rect 76076 84914 76132 84926
rect 77308 84308 77364 86382
rect 77868 86100 77924 86606
rect 78092 86436 78148 86446
rect 77868 86034 77924 86044
rect 77980 86434 78148 86436
rect 77980 86382 78094 86434
rect 78146 86382 78148 86434
rect 77980 86380 78148 86382
rect 77420 85764 77476 85774
rect 77420 85670 77476 85708
rect 77980 84420 78036 86380
rect 78092 86370 78148 86380
rect 78204 85986 78260 85998
rect 78204 85934 78206 85986
rect 78258 85934 78260 85986
rect 78204 85764 78260 85934
rect 78204 85698 78260 85708
rect 78092 84420 78148 84430
rect 77980 84418 78148 84420
rect 77980 84366 78094 84418
rect 78146 84366 78148 84418
rect 77980 84364 78148 84366
rect 78092 84354 78148 84364
rect 77420 84308 77476 84318
rect 77308 84252 77420 84308
rect 77420 84214 77476 84252
rect 76412 84194 76468 84206
rect 76412 84142 76414 84194
rect 76466 84142 76468 84194
rect 76412 84084 76468 84142
rect 76412 84018 76468 84028
rect 77420 84084 77476 84094
rect 76412 83412 76468 83422
rect 76412 83318 76468 83356
rect 77420 83410 77476 84028
rect 77420 83358 77422 83410
rect 77474 83358 77476 83410
rect 77420 83346 77476 83358
rect 77532 83522 77588 83534
rect 77532 83470 77534 83522
rect 77586 83470 77588 83522
rect 76076 83298 76132 83310
rect 76076 83246 76078 83298
rect 76130 83246 76132 83298
rect 76076 82852 76132 83246
rect 76188 82852 76244 82862
rect 76076 82850 76244 82852
rect 76076 82798 76190 82850
rect 76242 82798 76244 82850
rect 76076 82796 76244 82798
rect 76188 82786 76244 82796
rect 77532 82292 77588 83470
rect 78204 83524 78260 83534
rect 78204 83522 78372 83524
rect 78204 83470 78206 83522
rect 78258 83470 78372 83522
rect 78204 83468 78372 83470
rect 78204 83458 78260 83468
rect 77532 82068 77588 82236
rect 78316 82626 78372 83468
rect 78316 82574 78318 82626
rect 78370 82574 78372 82626
rect 77532 82002 77588 82012
rect 77868 82068 77924 82078
rect 77868 81974 77924 82012
rect 75740 81666 75796 81676
rect 76524 81732 76580 81742
rect 76524 81638 76580 81676
rect 77196 81732 77252 81742
rect 77308 81732 77364 81742
rect 77252 81730 77364 81732
rect 77252 81678 77310 81730
rect 77362 81678 77364 81730
rect 77252 81676 77364 81678
rect 75180 81564 75460 81620
rect 75068 81396 75124 81406
rect 75068 81302 75124 81340
rect 75292 81396 75348 81406
rect 74844 81116 75124 81172
rect 74396 80276 74452 80668
rect 74732 80658 74788 80668
rect 74508 80500 74564 80510
rect 74508 80406 74564 80444
rect 74956 80276 75012 80286
rect 74396 80274 75012 80276
rect 74396 80222 74958 80274
rect 75010 80222 75012 80274
rect 74396 80220 75012 80222
rect 74172 79714 74340 79716
rect 74172 79662 74174 79714
rect 74226 79662 74340 79714
rect 74172 79660 74340 79662
rect 74172 79650 74228 79660
rect 73836 78878 73838 78930
rect 73890 78878 73892 78930
rect 73836 78866 73892 78878
rect 74172 78708 74228 78718
rect 73948 78036 74004 78046
rect 73500 78034 74004 78036
rect 73500 77982 73950 78034
rect 74002 77982 74004 78034
rect 73500 77980 74004 77982
rect 73164 77924 73220 77934
rect 73276 77924 73332 77934
rect 73220 77922 73332 77924
rect 73220 77870 73278 77922
rect 73330 77870 73332 77922
rect 73220 77868 73332 77870
rect 72828 77422 72830 77474
rect 72882 77422 72884 77474
rect 72828 77410 72884 77422
rect 72940 77812 72996 77822
rect 72156 77140 72212 77150
rect 72156 77046 72212 77084
rect 72716 77140 72772 77150
rect 72716 77046 72772 77084
rect 72828 77140 72884 77150
rect 72940 77140 72996 77756
rect 72828 77138 72996 77140
rect 72828 77086 72830 77138
rect 72882 77086 72996 77138
rect 72828 77084 72996 77086
rect 72828 77074 72884 77084
rect 72156 76916 72212 76926
rect 72156 76354 72212 76860
rect 72156 76302 72158 76354
rect 72210 76302 72212 76354
rect 72156 76132 72212 76302
rect 72604 76356 72660 76366
rect 72604 76262 72660 76300
rect 72156 76066 72212 76076
rect 72828 76244 72884 76254
rect 72044 75730 72100 75740
rect 71932 75684 71988 75694
rect 71484 75012 71540 75022
rect 71036 75010 71540 75012
rect 71036 74958 71486 75010
rect 71538 74958 71540 75010
rect 71036 74956 71540 74958
rect 70924 74898 71428 74900
rect 70924 74846 70926 74898
rect 70978 74846 71428 74898
rect 70924 74844 71428 74846
rect 70924 74834 70980 74844
rect 69916 74788 69972 74798
rect 69804 74786 69972 74788
rect 69804 74734 69918 74786
rect 69970 74734 69972 74786
rect 69804 74732 69972 74734
rect 69804 74114 69860 74732
rect 69916 74722 69972 74732
rect 69804 74062 69806 74114
rect 69858 74062 69860 74114
rect 69804 73220 69860 74062
rect 70028 74002 70084 74014
rect 70028 73950 70030 74002
rect 70082 73950 70084 74002
rect 70028 73892 70084 73950
rect 70588 74004 70644 74014
rect 70588 73910 70644 73948
rect 70028 73826 70084 73836
rect 71260 73892 71316 73902
rect 71260 73798 71316 73836
rect 69804 73154 69860 73164
rect 71148 73220 71204 73230
rect 70812 72436 70868 72446
rect 70812 72342 70868 72380
rect 70476 72324 70532 72334
rect 69244 72322 69636 72324
rect 69244 72270 69246 72322
rect 69298 72270 69636 72322
rect 69244 72268 69636 72270
rect 70252 72322 70532 72324
rect 70252 72270 70478 72322
rect 70530 72270 70532 72322
rect 70252 72268 70532 72270
rect 69244 72258 69300 72268
rect 68908 71874 68964 71886
rect 68908 71822 68910 71874
rect 68962 71822 68964 71874
rect 68684 71762 68740 71774
rect 68684 71710 68686 71762
rect 68738 71710 68740 71762
rect 68572 70868 68628 70878
rect 68572 70774 68628 70812
rect 68684 69636 68740 71710
rect 68684 69570 68740 69580
rect 68796 70756 68852 70766
rect 68572 69300 68628 69310
rect 68572 69298 68740 69300
rect 68572 69246 68574 69298
rect 68626 69246 68740 69298
rect 68572 69244 68740 69246
rect 68572 69234 68628 69244
rect 68348 68226 68404 68236
rect 68460 69186 68516 69198
rect 68460 69134 68462 69186
rect 68514 69134 68516 69186
rect 68460 68068 68516 69134
rect 67676 68012 67844 68068
rect 67900 68066 68516 68068
rect 67900 68014 68462 68066
rect 68514 68014 68516 68066
rect 67900 68012 68516 68014
rect 67676 67730 67732 68012
rect 67788 67844 67844 67854
rect 67900 67844 67956 68012
rect 68460 68002 68516 68012
rect 67788 67842 67956 67844
rect 67788 67790 67790 67842
rect 67842 67790 67956 67842
rect 67788 67788 67956 67790
rect 67788 67778 67844 67788
rect 67676 67678 67678 67730
rect 67730 67678 67732 67730
rect 67676 67666 67732 67678
rect 68460 67732 68516 67742
rect 68460 67638 68516 67676
rect 68572 67730 68628 67742
rect 68572 67678 68574 67730
rect 68626 67678 68628 67730
rect 67564 67554 67620 67564
rect 68572 67508 68628 67678
rect 68572 67442 68628 67452
rect 68684 67396 68740 69244
rect 68684 67330 68740 67340
rect 68796 67172 68852 70700
rect 68908 70306 68964 71822
rect 69356 70978 69412 72268
rect 70252 71874 70308 72268
rect 70476 72258 70532 72268
rect 70252 71822 70254 71874
rect 70306 71822 70308 71874
rect 70252 71810 70308 71822
rect 69580 71762 69636 71774
rect 69580 71710 69582 71762
rect 69634 71710 69636 71762
rect 69580 71092 69636 71710
rect 69580 71026 69636 71036
rect 69356 70926 69358 70978
rect 69410 70926 69412 70978
rect 68908 70254 68910 70306
rect 68962 70254 68964 70306
rect 68908 70242 68964 70254
rect 69132 70532 69188 70542
rect 69020 68514 69076 68526
rect 69020 68462 69022 68514
rect 69074 68462 69076 68514
rect 69020 67732 69076 68462
rect 69132 67956 69188 70476
rect 69244 69524 69300 69534
rect 69244 69430 69300 69468
rect 69356 69412 69412 70926
rect 71036 70084 71092 70094
rect 70252 69636 70308 69646
rect 70252 69542 70308 69580
rect 69356 69346 69412 69356
rect 70588 69412 70644 69422
rect 71036 69412 71092 70028
rect 70588 69410 71092 69412
rect 70588 69358 70590 69410
rect 70642 69358 71092 69410
rect 70588 69356 71092 69358
rect 70588 68852 70644 69356
rect 70588 68786 70644 68796
rect 69580 68514 69636 68526
rect 69580 68462 69582 68514
rect 69634 68462 69636 68514
rect 69580 68404 69636 68462
rect 69916 68516 69972 68526
rect 69916 68422 69972 68460
rect 70588 68516 70644 68526
rect 71036 68516 71092 68526
rect 70588 68514 70756 68516
rect 70588 68462 70590 68514
rect 70642 68462 70756 68514
rect 70588 68460 70756 68462
rect 70588 68450 70644 68460
rect 69244 67956 69300 67966
rect 69132 67954 69412 67956
rect 69132 67902 69246 67954
rect 69298 67902 69412 67954
rect 69132 67900 69412 67902
rect 69244 67890 69300 67900
rect 69020 67666 69076 67676
rect 67340 67118 67342 67170
rect 67394 67118 67396 67170
rect 67340 67106 67396 67118
rect 68684 67116 68852 67172
rect 67452 66948 67508 66958
rect 67340 64932 67396 64942
rect 67340 64708 67396 64876
rect 67340 64642 67396 64652
rect 67340 64372 67396 64382
rect 67340 63924 67396 64316
rect 67340 63028 67396 63868
rect 67452 63922 67508 66892
rect 67788 66836 67844 66846
rect 67788 66386 67844 66780
rect 67788 66334 67790 66386
rect 67842 66334 67844 66386
rect 67788 66322 67844 66334
rect 67452 63870 67454 63922
rect 67506 63870 67508 63922
rect 67452 63858 67508 63870
rect 67564 66274 67620 66286
rect 67564 66222 67566 66274
rect 67618 66222 67620 66274
rect 67452 63028 67508 63038
rect 67340 63026 67508 63028
rect 67340 62974 67454 63026
rect 67506 62974 67508 63026
rect 67340 62972 67508 62974
rect 67452 62962 67508 62972
rect 67564 61684 67620 66222
rect 68572 66276 68628 66286
rect 68572 66182 68628 66220
rect 67900 66164 67956 66174
rect 67900 66070 67956 66108
rect 67676 66050 67732 66062
rect 67676 65998 67678 66050
rect 67730 65998 67732 66050
rect 67676 64708 67732 65998
rect 68012 66050 68068 66062
rect 68012 65998 68014 66050
rect 68066 65998 68068 66050
rect 67788 65156 67844 65166
rect 67788 64818 67844 65100
rect 67788 64766 67790 64818
rect 67842 64766 67844 64818
rect 67788 64754 67844 64766
rect 67676 64642 67732 64652
rect 67676 64036 67732 64046
rect 67676 64034 67956 64036
rect 67676 63982 67678 64034
rect 67730 63982 67956 64034
rect 67676 63980 67956 63982
rect 67676 63970 67732 63980
rect 67900 63138 67956 63980
rect 68012 63252 68068 65998
rect 68348 65380 68404 65390
rect 68124 64932 68180 64942
rect 68124 64818 68180 64876
rect 68124 64766 68126 64818
rect 68178 64766 68180 64818
rect 68124 64754 68180 64766
rect 68236 64596 68292 64606
rect 68124 63252 68180 63262
rect 68012 63250 68180 63252
rect 68012 63198 68126 63250
rect 68178 63198 68180 63250
rect 68012 63196 68180 63198
rect 68124 63186 68180 63196
rect 67900 63086 67902 63138
rect 67954 63086 67956 63138
rect 67900 63074 67956 63086
rect 68236 63138 68292 64540
rect 68348 63924 68404 65324
rect 68348 63792 68404 63868
rect 68460 64932 68516 64942
rect 68236 63086 68238 63138
rect 68290 63086 68292 63138
rect 68236 63074 68292 63086
rect 68460 63138 68516 64876
rect 68572 64596 68628 64606
rect 68572 64502 68628 64540
rect 68460 63086 68462 63138
rect 68514 63086 68516 63138
rect 68460 63074 68516 63086
rect 68684 62188 68740 67116
rect 68796 66836 68852 66846
rect 68796 63922 68852 66780
rect 69356 66274 69412 67900
rect 69580 67508 69636 68348
rect 70588 68292 70644 68302
rect 69916 67620 69972 67630
rect 69580 67442 69636 67452
rect 69804 67618 69972 67620
rect 69804 67566 69918 67618
rect 69970 67566 69972 67618
rect 69804 67564 69972 67566
rect 69468 66948 69524 66958
rect 69468 66854 69524 66892
rect 69356 66222 69358 66274
rect 69410 66222 69412 66274
rect 69356 66210 69412 66222
rect 69804 66276 69860 67564
rect 69916 67554 69972 67564
rect 70588 67618 70644 68236
rect 70588 67566 70590 67618
rect 70642 67566 70644 67618
rect 69916 67396 69972 67406
rect 69916 67170 69972 67340
rect 69916 67118 69918 67170
rect 69970 67118 69972 67170
rect 69916 67106 69972 67118
rect 70140 67170 70196 67182
rect 70140 67118 70142 67170
rect 70194 67118 70196 67170
rect 70140 66948 70196 67118
rect 70252 67172 70308 67182
rect 70252 67078 70308 67116
rect 70140 66882 70196 66892
rect 69692 66164 69748 66174
rect 69692 66070 69748 66108
rect 69468 66050 69524 66062
rect 69468 65998 69470 66050
rect 69522 65998 69524 66050
rect 69468 65940 69524 65998
rect 69468 65874 69524 65884
rect 69804 65940 69860 66220
rect 70476 66052 70532 66062
rect 69804 65874 69860 65884
rect 70364 66050 70532 66052
rect 70364 65998 70478 66050
rect 70530 65998 70532 66050
rect 70364 65996 70532 65998
rect 69244 65716 69300 65726
rect 69244 65490 69300 65660
rect 69244 65438 69246 65490
rect 69298 65438 69300 65490
rect 69244 65426 69300 65438
rect 69692 65156 69748 65166
rect 69692 64706 69748 65100
rect 70364 65044 70420 65996
rect 70476 65986 70532 65996
rect 69692 64654 69694 64706
rect 69746 64654 69748 64706
rect 69692 64642 69748 64654
rect 70140 64988 70364 65044
rect 69356 64596 69412 64606
rect 69356 64502 69412 64540
rect 68796 63870 68798 63922
rect 68850 63870 68852 63922
rect 68796 63858 68852 63870
rect 68908 64260 68964 64270
rect 68908 62804 68964 64204
rect 69692 63924 69748 63934
rect 69468 63922 69748 63924
rect 69468 63870 69694 63922
rect 69746 63870 69748 63922
rect 69468 63868 69748 63870
rect 69244 63028 69300 63038
rect 69244 62934 69300 62972
rect 68908 62738 68964 62748
rect 69244 62242 69300 62254
rect 69244 62190 69246 62242
rect 69298 62190 69300 62242
rect 69244 62188 69300 62190
rect 69468 62188 69524 63868
rect 69692 63858 69748 63868
rect 70140 63140 70196 64988
rect 70364 64978 70420 64988
rect 70476 64932 70532 64942
rect 70476 64594 70532 64876
rect 70476 64542 70478 64594
rect 70530 64542 70532 64594
rect 70476 64530 70532 64542
rect 70588 64372 70644 67566
rect 70700 67172 70756 68460
rect 70700 67106 70756 67116
rect 70924 68514 71092 68516
rect 70924 68462 71038 68514
rect 71090 68462 71092 68514
rect 70924 68460 71092 68462
rect 70700 66946 70756 66958
rect 70700 66894 70702 66946
rect 70754 66894 70756 66946
rect 70700 65604 70756 66894
rect 70924 66388 70980 68460
rect 71036 68450 71092 68460
rect 71148 68292 71204 73164
rect 71372 71316 71428 74844
rect 71484 74004 71540 74956
rect 71708 74898 71764 74910
rect 71708 74846 71710 74898
rect 71762 74846 71764 74898
rect 71708 74676 71764 74846
rect 71708 74610 71764 74620
rect 71484 73938 71540 73948
rect 71932 74002 71988 75628
rect 72268 74786 72324 74798
rect 72268 74734 72270 74786
rect 72322 74734 72324 74786
rect 72268 74676 72324 74734
rect 72268 74610 72324 74620
rect 71932 73950 71934 74002
rect 71986 73950 71988 74002
rect 71932 73938 71988 73950
rect 72268 74004 72324 74014
rect 72268 73910 72324 73948
rect 72716 74004 72772 74014
rect 72716 73910 72772 73948
rect 71708 73892 71764 73902
rect 71708 72658 71764 73836
rect 72492 73220 72548 73230
rect 71708 72606 71710 72658
rect 71762 72606 71764 72658
rect 71708 72594 71764 72606
rect 72268 73218 72548 73220
rect 72268 73166 72494 73218
rect 72546 73166 72548 73218
rect 72268 73164 72548 73166
rect 72268 72546 72324 73164
rect 72492 73154 72548 73164
rect 72828 72548 72884 76188
rect 72268 72494 72270 72546
rect 72322 72494 72324 72546
rect 72156 72436 72212 72446
rect 72044 71652 72100 71662
rect 71372 71260 71540 71316
rect 71372 71092 71428 71102
rect 71372 70998 71428 71036
rect 71484 70868 71540 71260
rect 71372 70644 71428 70654
rect 71372 69748 71428 70588
rect 71260 69692 71428 69748
rect 71484 70418 71540 70812
rect 71484 70366 71486 70418
rect 71538 70366 71540 70418
rect 71260 69410 71316 69692
rect 71484 69636 71540 70366
rect 72044 70644 72100 71596
rect 72044 70194 72100 70588
rect 72044 70142 72046 70194
rect 72098 70142 72100 70194
rect 72044 70130 72100 70142
rect 71484 69570 71540 69580
rect 72156 69634 72212 72380
rect 72268 72100 72324 72494
rect 72268 72034 72324 72044
rect 72716 72492 72884 72548
rect 72604 71988 72660 71998
rect 72156 69582 72158 69634
rect 72210 69582 72212 69634
rect 72156 69570 72212 69582
rect 72380 71650 72436 71662
rect 72380 71598 72382 71650
rect 72434 71598 72436 71650
rect 71260 69358 71262 69410
rect 71314 69358 71316 69410
rect 71260 69346 71316 69358
rect 71372 69300 71428 69310
rect 71372 69206 71428 69244
rect 72380 69300 72436 71598
rect 72604 70418 72660 71932
rect 72604 70366 72606 70418
rect 72658 70366 72660 70418
rect 72604 70354 72660 70366
rect 72716 69972 72772 72492
rect 72828 72322 72884 72334
rect 72828 72270 72830 72322
rect 72882 72270 72884 72322
rect 72828 70084 72884 72270
rect 72828 70018 72884 70028
rect 72604 69916 72772 69972
rect 72492 69636 72548 69646
rect 72492 69542 72548 69580
rect 72380 69234 72436 69244
rect 71036 68236 71204 68292
rect 71372 68514 71428 68526
rect 71372 68462 71374 68514
rect 71426 68462 71428 68514
rect 71036 66948 71092 68236
rect 71372 68180 71428 68462
rect 71372 68114 71428 68124
rect 71820 68516 71876 68526
rect 71148 67620 71204 67630
rect 71596 67620 71652 67630
rect 71148 67618 71540 67620
rect 71148 67566 71150 67618
rect 71202 67566 71540 67618
rect 71148 67564 71540 67566
rect 71148 67554 71204 67564
rect 71148 66948 71204 66958
rect 71036 66946 71204 66948
rect 71036 66894 71150 66946
rect 71202 66894 71204 66946
rect 71036 66892 71204 66894
rect 71148 66836 71204 66892
rect 71148 66770 71204 66780
rect 70924 66332 71092 66388
rect 70700 65538 70756 65548
rect 70812 66164 70868 66174
rect 70812 65380 70868 66108
rect 70924 66050 70980 66062
rect 70924 65998 70926 66050
rect 70978 65998 70980 66050
rect 70924 65828 70980 65998
rect 71036 66052 71092 66332
rect 71036 65986 71092 65996
rect 71260 66050 71316 66062
rect 71260 65998 71262 66050
rect 71314 65998 71316 66050
rect 70924 65762 70980 65772
rect 71148 65492 71204 65502
rect 71148 65398 71204 65436
rect 70700 65324 70868 65380
rect 70700 64484 70756 65324
rect 70924 65266 70980 65278
rect 70924 65214 70926 65266
rect 70978 65214 70980 65266
rect 70812 64708 70868 64718
rect 70924 64708 70980 65214
rect 71260 64932 71316 65998
rect 71484 65492 71540 67564
rect 71596 67526 71652 67564
rect 71820 67282 71876 68460
rect 71820 67230 71822 67282
rect 71874 67230 71876 67282
rect 71820 67218 71876 67230
rect 71932 68514 71988 68526
rect 71932 68462 71934 68514
rect 71986 68462 71988 68514
rect 71932 66724 71988 68462
rect 72492 68514 72548 68526
rect 72492 68462 72494 68514
rect 72546 68462 72548 68514
rect 72492 68292 72548 68462
rect 72492 68226 72548 68236
rect 72604 67954 72660 69916
rect 73052 69300 73108 69310
rect 73052 69206 73108 69244
rect 72604 67902 72606 67954
rect 72658 67902 72660 67954
rect 72604 67890 72660 67902
rect 72492 67842 72548 67854
rect 72492 67790 72494 67842
rect 72546 67790 72548 67842
rect 72044 67620 72100 67630
rect 72044 67526 72100 67564
rect 72268 67620 72324 67630
rect 72156 67058 72212 67070
rect 72156 67006 72158 67058
rect 72210 67006 72212 67058
rect 72156 66948 72212 67006
rect 72156 66882 72212 66892
rect 71932 66612 71988 66668
rect 71820 66556 71988 66612
rect 71708 66050 71764 66062
rect 71708 65998 71710 66050
rect 71762 65998 71764 66050
rect 71596 65492 71652 65502
rect 71484 65490 71652 65492
rect 71484 65438 71598 65490
rect 71650 65438 71652 65490
rect 71484 65436 71652 65438
rect 71484 65266 71540 65436
rect 71596 65426 71652 65436
rect 71484 65214 71486 65266
rect 71538 65214 71540 65266
rect 71484 65202 71540 65214
rect 71708 65266 71764 65998
rect 71708 65214 71710 65266
rect 71762 65214 71764 65266
rect 71708 65202 71764 65214
rect 71820 64932 71876 66556
rect 72044 65380 72100 65390
rect 72044 65286 72100 65324
rect 71260 64866 71316 64876
rect 71484 64876 71876 64932
rect 71932 65266 71988 65278
rect 71932 65214 71934 65266
rect 71986 65214 71988 65266
rect 70812 64706 70980 64708
rect 70812 64654 70814 64706
rect 70866 64654 70980 64706
rect 70812 64652 70980 64654
rect 70812 64642 70868 64652
rect 70700 64428 70868 64484
rect 70588 64316 70756 64372
rect 70588 64036 70644 64046
rect 70588 63588 70644 63980
rect 70700 63700 70756 64316
rect 70700 63634 70756 63644
rect 70476 63532 70644 63588
rect 70140 63138 70420 63140
rect 70140 63086 70142 63138
rect 70194 63086 70420 63138
rect 70140 63084 70420 63086
rect 70140 63074 70196 63084
rect 69916 63028 69972 63038
rect 69804 62916 69860 62926
rect 68684 62132 68852 62188
rect 69244 62132 69524 62188
rect 69692 62914 69860 62916
rect 69692 62862 69806 62914
rect 69858 62862 69860 62914
rect 69692 62860 69860 62862
rect 67900 61684 67956 61694
rect 67564 61682 67956 61684
rect 67564 61630 67902 61682
rect 67954 61630 67956 61682
rect 67564 61628 67956 61630
rect 67900 61618 67956 61628
rect 68236 61684 68292 61694
rect 67452 61572 67508 61582
rect 67452 61478 67508 61516
rect 68124 61570 68180 61582
rect 68124 61518 68126 61570
rect 68178 61518 68180 61570
rect 67676 61460 67732 61470
rect 67676 61366 67732 61404
rect 67228 61292 67508 61348
rect 67228 60900 67284 60910
rect 67228 60898 67396 60900
rect 67228 60846 67230 60898
rect 67282 60846 67396 60898
rect 67228 60844 67396 60846
rect 67228 60834 67284 60844
rect 67116 60722 67172 60732
rect 66892 60508 67172 60564
rect 66780 60174 66782 60226
rect 66834 60174 66836 60226
rect 66780 60162 66836 60174
rect 66780 59892 66836 59902
rect 66780 59798 66836 59836
rect 66668 59612 67060 59668
rect 66556 59276 66836 59332
rect 66444 59164 66612 59220
rect 65884 59154 65940 59164
rect 65772 59108 65828 59118
rect 65772 58322 65828 59052
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65772 58270 65774 58322
rect 65826 58270 65828 58322
rect 65772 58258 65828 58270
rect 65884 58436 65940 58446
rect 65884 58322 65940 58380
rect 65884 58270 65886 58322
rect 65938 58270 65940 58322
rect 65660 58146 65716 58156
rect 65884 58212 65940 58270
rect 66108 58212 66164 58222
rect 65884 58156 66108 58212
rect 65324 57822 65326 57874
rect 65378 57822 65380 57874
rect 65324 57810 65380 57822
rect 65548 57876 65604 57886
rect 65548 57782 65604 57820
rect 65660 57764 65716 57774
rect 65884 57764 65940 58156
rect 66108 57874 66164 58156
rect 66444 58212 66500 58222
rect 66444 58118 66500 58156
rect 66108 57822 66110 57874
rect 66162 57822 66164 57874
rect 66108 57810 66164 57822
rect 65660 57762 65940 57764
rect 65660 57710 65662 57762
rect 65714 57710 65940 57762
rect 65660 57708 65940 57710
rect 65660 57698 65716 57708
rect 64764 57538 64820 57550
rect 64764 57486 64766 57538
rect 64818 57486 64820 57538
rect 64764 57092 64820 57486
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 64764 57026 64820 57036
rect 64764 56644 64820 56654
rect 65212 56644 65268 56654
rect 64764 56642 65268 56644
rect 64764 56590 64766 56642
rect 64818 56590 65214 56642
rect 65266 56590 65268 56642
rect 64764 56588 65268 56590
rect 64764 55188 64820 56588
rect 65212 56578 65268 56588
rect 65548 56196 65604 56206
rect 65548 56102 65604 56140
rect 64764 55122 64820 55132
rect 65324 56082 65380 56094
rect 65324 56030 65326 56082
rect 65378 56030 65380 56082
rect 65324 55076 65380 56030
rect 65660 56084 65716 56094
rect 66108 56084 66164 56094
rect 65660 56082 66164 56084
rect 65660 56030 65662 56082
rect 65714 56030 66110 56082
rect 66162 56030 66164 56082
rect 65660 56028 66164 56030
rect 65660 55468 65716 56028
rect 66108 56018 66164 56028
rect 66444 55860 66500 55870
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 65324 55010 65380 55020
rect 65548 55412 65716 55468
rect 65324 54740 65380 54750
rect 64764 53732 64820 53742
rect 64652 53730 64820 53732
rect 64652 53678 64766 53730
rect 64818 53678 64820 53730
rect 64652 53676 64820 53678
rect 64764 53666 64820 53676
rect 65324 53730 65380 54684
rect 65548 54180 65604 55412
rect 65660 55188 65716 55198
rect 65660 54516 65716 55132
rect 66444 54626 66500 55804
rect 66556 55468 66612 59164
rect 66780 55468 66836 59276
rect 66892 59218 66948 59230
rect 66892 59166 66894 59218
rect 66946 59166 66948 59218
rect 66892 59108 66948 59166
rect 66892 59042 66948 59052
rect 67004 58548 67060 59612
rect 66892 58212 66948 58222
rect 66892 56756 66948 58156
rect 67004 57650 67060 58492
rect 67004 57598 67006 57650
rect 67058 57598 67060 57650
rect 67004 57586 67060 57598
rect 66892 56690 66948 56700
rect 67116 56644 67172 60508
rect 67228 60116 67284 60126
rect 67228 60022 67284 60060
rect 67340 60004 67396 60844
rect 67452 60788 67508 61292
rect 67564 60788 67620 60798
rect 67452 60786 67620 60788
rect 67452 60734 67566 60786
rect 67618 60734 67620 60786
rect 67452 60732 67620 60734
rect 67564 60452 67620 60732
rect 67564 60386 67620 60396
rect 67676 60788 67732 60798
rect 67340 59218 67396 59948
rect 67676 60002 67732 60732
rect 67676 59950 67678 60002
rect 67730 59950 67732 60002
rect 67676 59938 67732 59950
rect 68012 60564 68068 60574
rect 68012 60002 68068 60508
rect 68012 59950 68014 60002
rect 68066 59950 68068 60002
rect 68012 59938 68068 59950
rect 67900 59780 67956 59790
rect 67340 59166 67342 59218
rect 67394 59166 67396 59218
rect 67340 59154 67396 59166
rect 67452 59778 67956 59780
rect 67452 59726 67902 59778
rect 67954 59726 67956 59778
rect 67452 59724 67956 59726
rect 67116 56578 67172 56588
rect 67452 56420 67508 59724
rect 67900 59714 67956 59724
rect 68124 59556 68180 61518
rect 68236 60898 68292 61628
rect 68460 61684 68516 61694
rect 68460 61590 68516 61628
rect 68796 61348 68852 62132
rect 69244 61796 69300 61806
rect 69244 61682 69300 61740
rect 69244 61630 69246 61682
rect 69298 61630 69300 61682
rect 69244 61460 69300 61630
rect 69244 61394 69300 61404
rect 68684 61292 68852 61348
rect 68236 60846 68238 60898
rect 68290 60846 68292 60898
rect 68236 60834 68292 60846
rect 68572 60898 68628 60910
rect 68572 60846 68574 60898
rect 68626 60846 68628 60898
rect 68460 60452 68516 60462
rect 68460 60114 68516 60396
rect 68460 60062 68462 60114
rect 68514 60062 68516 60114
rect 68460 60050 68516 60062
rect 68572 60004 68628 60846
rect 68572 59938 68628 59948
rect 68572 59780 68628 59790
rect 67900 59500 68180 59556
rect 68460 59556 68516 59566
rect 67900 59442 67956 59500
rect 67900 59390 67902 59442
rect 67954 59390 67956 59442
rect 67900 59378 67956 59390
rect 68124 59218 68180 59230
rect 68124 59166 68126 59218
rect 68178 59166 68180 59218
rect 68124 58548 68180 59166
rect 68124 58482 68180 58492
rect 68236 58436 68292 58446
rect 68236 58342 68292 58380
rect 67564 57650 67620 57662
rect 67564 57598 67566 57650
rect 67618 57598 67620 57650
rect 67564 57540 67620 57598
rect 68012 57540 68068 57550
rect 68124 57540 68180 57550
rect 67564 57538 68124 57540
rect 67564 57486 68014 57538
rect 68066 57486 68124 57538
rect 67564 57484 68124 57486
rect 68012 57474 68068 57484
rect 68124 56866 68180 57484
rect 68124 56814 68126 56866
rect 68178 56814 68180 56866
rect 67452 56364 67620 56420
rect 67564 56308 67620 56364
rect 68012 56308 68068 56318
rect 67564 56306 68068 56308
rect 67564 56254 68014 56306
rect 68066 56254 68068 56306
rect 67564 56252 68068 56254
rect 67452 56196 67508 56206
rect 67340 56194 67508 56196
rect 67340 56142 67454 56194
rect 67506 56142 67508 56194
rect 67340 56140 67508 56142
rect 66556 55412 66724 55468
rect 66780 55412 66948 55468
rect 66444 54574 66446 54626
rect 66498 54574 66500 54626
rect 66444 54562 66500 54574
rect 65660 54514 65828 54516
rect 65660 54462 65662 54514
rect 65714 54462 65828 54514
rect 65660 54460 65828 54462
rect 65660 54450 65716 54460
rect 65548 54124 65716 54180
rect 65324 53678 65326 53730
rect 65378 53678 65380 53730
rect 65324 53666 65380 53678
rect 65548 53844 65604 53854
rect 64540 53620 64596 53630
rect 64540 53060 64596 53564
rect 65548 53618 65604 53788
rect 65548 53566 65550 53618
rect 65602 53566 65604 53618
rect 65548 53554 65604 53566
rect 65660 53620 65716 54124
rect 65660 53526 65716 53564
rect 65324 53172 65380 53182
rect 65772 53172 65828 54460
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 66108 53620 66164 53630
rect 66108 53526 66164 53564
rect 65324 53170 66612 53172
rect 65324 53118 65326 53170
rect 65378 53118 65774 53170
rect 65826 53118 66612 53170
rect 65324 53116 66612 53118
rect 65324 53106 65380 53116
rect 65772 53106 65828 53116
rect 64540 52966 64596 53004
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 66332 52274 66388 53116
rect 66556 52946 66612 53116
rect 66556 52894 66558 52946
rect 66610 52894 66612 52946
rect 66556 52882 66612 52894
rect 66332 52222 66334 52274
rect 66386 52222 66388 52274
rect 66332 52210 66388 52222
rect 64764 51604 64820 51614
rect 64540 51380 64596 51390
rect 64540 51266 64596 51324
rect 64540 51214 64542 51266
rect 64594 51214 64596 51266
rect 64540 50484 64596 51214
rect 64764 50706 64820 51548
rect 65324 51604 65380 51614
rect 65324 51510 65380 51548
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 64764 50654 64766 50706
rect 64818 50654 64820 50706
rect 64764 50642 64820 50654
rect 65996 50818 66052 50830
rect 65996 50766 65998 50818
rect 66050 50766 66052 50818
rect 65996 50706 66052 50766
rect 66556 50820 66612 50830
rect 66668 50820 66724 55412
rect 66556 50818 66724 50820
rect 66556 50766 66558 50818
rect 66610 50766 66724 50818
rect 66556 50764 66724 50766
rect 66556 50754 66612 50764
rect 65996 50654 65998 50706
rect 66050 50654 66052 50706
rect 64540 50418 64596 50428
rect 65324 50484 65380 50494
rect 65324 50390 65380 50428
rect 65436 50372 65492 50382
rect 65324 49812 65380 49822
rect 65324 49718 65380 49756
rect 64652 49700 64708 49710
rect 64652 49606 64708 49644
rect 65436 49700 65492 50316
rect 65660 50370 65716 50382
rect 65660 50318 65662 50370
rect 65714 50318 65716 50370
rect 65436 49634 65492 49644
rect 65548 49922 65604 49934
rect 65548 49870 65550 49922
rect 65602 49870 65604 49922
rect 65548 49028 65604 49870
rect 65660 49922 65716 50318
rect 65996 50372 66052 50654
rect 65996 50306 66052 50316
rect 66444 50484 66500 50494
rect 66444 50370 66500 50428
rect 66892 50428 66948 55412
rect 67004 53732 67060 53742
rect 67340 53732 67396 56140
rect 67452 56130 67508 56140
rect 67564 56194 67620 56252
rect 68012 56242 68068 56252
rect 67564 56142 67566 56194
rect 67618 56142 67620 56194
rect 67564 56130 67620 56142
rect 67452 55860 67508 55870
rect 67452 55766 67508 55804
rect 68124 55412 68180 56814
rect 68460 56868 68516 59500
rect 68572 59332 68628 59724
rect 68572 59218 68628 59276
rect 68572 59166 68574 59218
rect 68626 59166 68628 59218
rect 68572 59154 68628 59166
rect 68572 58436 68628 58446
rect 68572 58342 68628 58380
rect 68572 56868 68628 56878
rect 68460 56866 68628 56868
rect 68460 56814 68574 56866
rect 68626 56814 68628 56866
rect 68460 56812 68628 56814
rect 68236 56308 68292 56318
rect 68236 56306 68516 56308
rect 68236 56254 68238 56306
rect 68290 56254 68516 56306
rect 68236 56252 68516 56254
rect 68236 56242 68292 56252
rect 68348 56084 68404 56094
rect 68348 55990 68404 56028
rect 68124 55346 68180 55356
rect 68460 54404 68516 56252
rect 68572 55748 68628 56812
rect 68572 55682 68628 55692
rect 68572 55298 68628 55310
rect 68572 55246 68574 55298
rect 68626 55246 68628 55298
rect 68572 55074 68628 55246
rect 68572 55022 68574 55074
rect 68626 55022 68628 55074
rect 68572 55010 68628 55022
rect 68572 54404 68628 54414
rect 68460 54402 68628 54404
rect 68460 54350 68574 54402
rect 68626 54350 68628 54402
rect 68460 54348 68628 54350
rect 68572 54338 68628 54348
rect 67452 53732 67508 53742
rect 67340 53730 67508 53732
rect 67340 53678 67454 53730
rect 67506 53678 67508 53730
rect 67340 53676 67508 53678
rect 67004 53638 67060 53676
rect 67452 53666 67508 53676
rect 67788 53732 67844 53742
rect 67788 53638 67844 53676
rect 68572 53618 68628 53630
rect 68572 53566 68574 53618
rect 68626 53566 68628 53618
rect 67676 53506 67732 53518
rect 67676 53454 67678 53506
rect 67730 53454 67732 53506
rect 67340 53060 67396 53070
rect 67340 52966 67396 53004
rect 67004 52612 67060 52622
rect 67004 52162 67060 52556
rect 67004 52110 67006 52162
rect 67058 52110 67060 52162
rect 67004 52098 67060 52110
rect 67116 52500 67172 52510
rect 67116 52050 67172 52444
rect 67676 52276 67732 53454
rect 68236 53506 68292 53518
rect 68236 53454 68238 53506
rect 68290 53454 68292 53506
rect 68236 53060 68292 53454
rect 68236 52994 68292 53004
rect 68460 53506 68516 53518
rect 68460 53454 68462 53506
rect 68514 53454 68516 53506
rect 68460 52276 68516 53454
rect 68572 53508 68628 53566
rect 68572 52500 68628 53452
rect 68572 52434 68628 52444
rect 67676 52220 67956 52276
rect 67116 51998 67118 52050
rect 67170 51998 67172 52050
rect 67116 51986 67172 51998
rect 67788 52052 67844 52062
rect 67788 51958 67844 51996
rect 67900 52050 67956 52220
rect 68124 52220 68516 52276
rect 68124 52162 68180 52220
rect 68572 52164 68628 52174
rect 68124 52110 68126 52162
rect 68178 52110 68180 52162
rect 68124 52098 68180 52110
rect 68460 52108 68572 52164
rect 67900 51998 67902 52050
rect 67954 51998 67956 52050
rect 67340 51940 67396 51950
rect 67340 51938 67732 51940
rect 67340 51886 67342 51938
rect 67394 51886 67732 51938
rect 67340 51884 67732 51886
rect 67340 51874 67396 51884
rect 67676 51716 67732 51884
rect 67900 51828 67956 51998
rect 68460 52050 68516 52108
rect 68572 52098 68628 52108
rect 68460 51998 68462 52050
rect 68514 51998 68516 52050
rect 68460 51986 68516 51998
rect 67900 51772 68404 51828
rect 67676 51660 68068 51716
rect 68012 51490 68068 51660
rect 68012 51438 68014 51490
rect 68066 51438 68068 51490
rect 68012 51426 68068 51438
rect 67340 51378 67396 51390
rect 67340 51326 67342 51378
rect 67394 51326 67396 51378
rect 67340 50596 67396 51326
rect 67340 50530 67396 50540
rect 66892 50372 67060 50428
rect 66444 50318 66446 50370
rect 66498 50318 66500 50370
rect 65660 49870 65662 49922
rect 65714 49870 65716 49922
rect 65660 49858 65716 49870
rect 66332 49924 66388 49934
rect 66332 49830 66388 49868
rect 66444 49810 66500 50318
rect 66444 49758 66446 49810
rect 66498 49758 66500 49810
rect 66332 49586 66388 49598
rect 66332 49534 66334 49586
rect 66386 49534 66388 49586
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65548 48972 65940 49028
rect 65212 48916 65268 48926
rect 65268 48860 65604 48916
rect 65212 48784 65268 48860
rect 65548 48804 65604 48860
rect 65548 48748 65828 48804
rect 65100 48580 65156 48590
rect 64988 47346 65044 47358
rect 64988 47294 64990 47346
rect 65042 47294 65044 47346
rect 64876 47236 64932 47246
rect 64876 45780 64932 47180
rect 64988 46114 65044 47294
rect 64988 46062 64990 46114
rect 65042 46062 65044 46114
rect 64988 46050 65044 46062
rect 65100 45890 65156 48524
rect 65548 48356 65604 48366
rect 65548 48262 65604 48300
rect 65100 45838 65102 45890
rect 65154 45838 65156 45890
rect 65100 45826 65156 45838
rect 65324 48242 65380 48254
rect 65324 48190 65326 48242
rect 65378 48190 65380 48242
rect 64988 45780 65044 45790
rect 64876 45778 65044 45780
rect 64876 45726 64990 45778
rect 65042 45726 65044 45778
rect 64876 45724 65044 45726
rect 64988 45714 65044 45724
rect 65324 45444 65380 48190
rect 65660 48242 65716 48254
rect 65660 48190 65662 48242
rect 65714 48190 65716 48242
rect 65436 48132 65492 48142
rect 65436 46452 65492 48076
rect 65660 47236 65716 48190
rect 65772 47458 65828 48748
rect 65884 48244 65940 48972
rect 66332 48580 66388 49534
rect 66444 49588 66500 49758
rect 66444 49522 66500 49532
rect 66892 49924 66948 49934
rect 66892 48692 66948 49868
rect 66892 48626 66948 48636
rect 66332 48514 66388 48524
rect 66332 48354 66388 48366
rect 67004 48356 67060 50372
rect 68348 50036 68404 51772
rect 68572 50596 68628 50606
rect 68348 50034 68516 50036
rect 68348 49982 68350 50034
rect 68402 49982 68516 50034
rect 68348 49980 68516 49982
rect 68348 49970 68404 49980
rect 68236 49924 68292 49934
rect 68012 49812 68068 49822
rect 67452 49698 67508 49710
rect 67452 49646 67454 49698
rect 67506 49646 67508 49698
rect 67452 49588 67508 49646
rect 67452 49522 67508 49532
rect 67116 49028 67172 49038
rect 67228 49028 67284 49038
rect 67116 49026 67228 49028
rect 67116 48974 67118 49026
rect 67170 48974 67228 49026
rect 67116 48972 67228 48974
rect 67116 48962 67172 48972
rect 66332 48302 66334 48354
rect 66386 48302 66388 48354
rect 65884 48178 65940 48188
rect 66108 48244 66164 48254
rect 66108 48150 66164 48188
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65772 47406 65774 47458
rect 65826 47406 65828 47458
rect 65772 47394 65828 47406
rect 66108 47460 66164 47470
rect 65660 47170 65716 47180
rect 66108 46900 66164 47404
rect 66220 47236 66276 47246
rect 66220 47142 66276 47180
rect 66332 47124 66388 48302
rect 66780 48300 67060 48356
rect 67116 48468 67172 48478
rect 66444 48244 66500 48254
rect 66444 48242 66612 48244
rect 66444 48190 66446 48242
rect 66498 48190 66612 48242
rect 66444 48188 66612 48190
rect 66444 48178 66500 48188
rect 66556 47460 66612 48188
rect 66556 47366 66612 47404
rect 66332 47058 66388 47068
rect 66444 47234 66500 47246
rect 66444 47182 66446 47234
rect 66498 47182 66500 47234
rect 66220 46900 66276 46910
rect 65660 46898 66276 46900
rect 65660 46846 66222 46898
rect 66274 46846 66276 46898
rect 65660 46844 66276 46846
rect 65548 46788 65604 46798
rect 65548 46694 65604 46732
rect 65660 46786 65716 46844
rect 66220 46834 66276 46844
rect 65660 46734 65662 46786
rect 65714 46734 65716 46786
rect 65660 46722 65716 46734
rect 65548 46452 65604 46462
rect 65436 46450 65604 46452
rect 65436 46398 65550 46450
rect 65602 46398 65604 46450
rect 65436 46396 65604 46398
rect 65548 46386 65604 46396
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65324 45378 65380 45388
rect 66444 44996 66500 47182
rect 66444 44930 66500 44940
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 64428 44492 64820 44548
rect 64204 43586 64260 43596
rect 64428 43650 64484 43662
rect 64428 43598 64430 43650
rect 64482 43598 64484 43650
rect 63756 43314 63812 43326
rect 63756 43262 63758 43314
rect 63810 43262 63812 43314
rect 63756 41972 63812 43262
rect 64428 43316 64484 43598
rect 64540 43540 64596 43550
rect 64540 43446 64596 43484
rect 64428 43250 64484 43260
rect 63868 42868 63924 42878
rect 63868 42774 63924 42812
rect 64316 42082 64372 42094
rect 64316 42030 64318 42082
rect 64370 42030 64372 42082
rect 63756 41916 64260 41972
rect 63420 41860 63476 41870
rect 63420 41766 63476 41804
rect 63756 41746 63812 41758
rect 63756 41694 63758 41746
rect 63810 41694 63812 41746
rect 63532 40516 63588 40526
rect 63532 40422 63588 40460
rect 63756 39396 63812 41694
rect 64204 41300 64260 41916
rect 64316 41748 64372 42030
rect 64316 41682 64372 41692
rect 64428 41970 64484 41982
rect 64428 41918 64430 41970
rect 64482 41918 64484 41970
rect 63980 40516 64036 40526
rect 63980 40422 64036 40460
rect 64204 40290 64260 41244
rect 64316 41524 64372 41534
rect 64316 41298 64372 41468
rect 64316 41246 64318 41298
rect 64370 41246 64372 41298
rect 64316 41234 64372 41246
rect 64428 41300 64484 41918
rect 64428 41234 64484 41244
rect 64652 41860 64708 41870
rect 64540 40628 64596 40638
rect 64652 40628 64708 41804
rect 64540 40626 64708 40628
rect 64540 40574 64542 40626
rect 64594 40574 64708 40626
rect 64540 40572 64708 40574
rect 64540 40562 64596 40572
rect 64204 40238 64206 40290
rect 64258 40238 64260 40290
rect 64204 40226 64260 40238
rect 63756 39330 63812 39340
rect 63980 38948 64036 38958
rect 63980 38854 64036 38892
rect 63420 38836 63476 38846
rect 63420 37490 63476 38780
rect 64204 38836 64260 38846
rect 64204 38742 64260 38780
rect 64764 38668 64820 44492
rect 66332 44210 66388 44222
rect 66332 44158 66334 44210
rect 66386 44158 66388 44210
rect 66332 43652 66388 44158
rect 65324 43540 65380 43550
rect 65324 43426 65380 43484
rect 65324 43374 65326 43426
rect 65378 43374 65380 43426
rect 64988 41188 65044 41198
rect 64988 39730 65044 41132
rect 64988 39678 64990 39730
rect 65042 39678 65044 39730
rect 64988 39666 65044 39678
rect 65212 40516 65268 40526
rect 65212 40404 65268 40460
rect 65324 40404 65380 43374
rect 65772 43540 65828 43550
rect 65772 43316 65828 43484
rect 65772 42980 65828 43260
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65772 42924 66052 42980
rect 65996 42866 66052 42924
rect 65996 42814 65998 42866
rect 66050 42814 66052 42866
rect 65996 42802 66052 42814
rect 65436 42082 65492 42094
rect 65436 42030 65438 42082
rect 65490 42030 65492 42082
rect 65436 41524 65492 42030
rect 65772 42084 65828 42094
rect 65772 41990 65828 42028
rect 66332 41970 66388 43596
rect 66780 43540 66836 48300
rect 66892 48132 66948 48170
rect 66892 48066 66948 48076
rect 66892 47908 66948 47918
rect 66892 46674 66948 47852
rect 67004 47572 67060 47582
rect 67116 47572 67172 48412
rect 67004 47570 67172 47572
rect 67004 47518 67006 47570
rect 67058 47518 67172 47570
rect 67004 47516 67172 47518
rect 67004 47460 67060 47516
rect 67004 47394 67060 47404
rect 66892 46622 66894 46674
rect 66946 46622 66948 46674
rect 66892 46610 66948 46622
rect 67004 45108 67060 45118
rect 67004 45014 67060 45052
rect 66780 43474 66836 43484
rect 67228 44322 67284 48972
rect 67452 48916 67508 48926
rect 67340 48468 67396 48478
rect 67340 48374 67396 48412
rect 67452 48132 67508 48860
rect 67452 48066 67508 48076
rect 67676 48804 67732 48814
rect 68012 48804 68068 49756
rect 68236 49028 68292 49868
rect 68348 49028 68404 49038
rect 68236 49026 68404 49028
rect 68236 48974 68350 49026
rect 68402 48974 68404 49026
rect 68236 48972 68404 48974
rect 68236 48916 68292 48972
rect 68348 48962 68404 48972
rect 68236 48850 68292 48860
rect 68460 48914 68516 49980
rect 68460 48862 68462 48914
rect 68514 48862 68516 48914
rect 67676 48802 68068 48804
rect 67676 48750 67678 48802
rect 67730 48750 68068 48802
rect 67676 48748 68068 48750
rect 67676 46900 67732 48748
rect 68460 48692 68516 48862
rect 68012 48636 68516 48692
rect 68012 48466 68068 48636
rect 68012 48414 68014 48466
rect 68066 48414 68068 48466
rect 68012 48402 68068 48414
rect 67900 48242 67956 48254
rect 67900 48190 67902 48242
rect 67954 48190 67956 48242
rect 67900 48020 67956 48190
rect 68236 48244 68292 48254
rect 68572 48244 68628 50540
rect 68684 49812 68740 61292
rect 69244 61012 69300 61022
rect 69356 61012 69412 62132
rect 69692 61572 69748 62860
rect 69804 62850 69860 62860
rect 69916 62354 69972 62972
rect 69916 62302 69918 62354
rect 69970 62302 69972 62354
rect 69916 62244 69972 62302
rect 70140 62356 70196 62366
rect 70140 62262 70196 62300
rect 69916 62178 69972 62188
rect 69692 61506 69748 61516
rect 70252 61572 70308 61582
rect 70252 61478 70308 61516
rect 70028 61460 70084 61470
rect 70028 61458 70196 61460
rect 70028 61406 70030 61458
rect 70082 61406 70196 61458
rect 70028 61404 70196 61406
rect 70028 61394 70084 61404
rect 69244 61010 69412 61012
rect 69244 60958 69246 61010
rect 69298 60958 69412 61010
rect 69244 60956 69412 60958
rect 70028 61236 70084 61246
rect 69244 60946 69300 60956
rect 69916 60900 69972 60910
rect 69356 60788 69412 60798
rect 69356 60694 69412 60732
rect 69244 60564 69300 60574
rect 69244 60470 69300 60508
rect 69804 60452 69860 60462
rect 69468 60004 69524 60014
rect 69356 59332 69412 59342
rect 69356 59238 69412 59276
rect 68908 59106 68964 59118
rect 68908 59054 68910 59106
rect 68962 59054 68964 59106
rect 68908 58660 68964 59054
rect 69244 59108 69300 59118
rect 69244 58772 69300 59052
rect 69244 58716 69412 58772
rect 69132 58660 69188 58670
rect 68908 58658 69188 58660
rect 68908 58606 69134 58658
rect 69186 58606 69188 58658
rect 68908 58604 69188 58606
rect 69132 58594 69188 58604
rect 69244 58548 69300 58558
rect 68796 57540 68852 57550
rect 68796 57446 68852 57484
rect 68908 56084 68964 56094
rect 68908 55990 68964 56028
rect 69244 55468 69300 58492
rect 69356 58546 69412 58716
rect 69356 58494 69358 58546
rect 69410 58494 69412 58546
rect 69356 58482 69412 58494
rect 69468 58324 69524 59948
rect 69804 59890 69860 60396
rect 69916 60116 69972 60844
rect 70028 60788 70084 61180
rect 70140 60900 70196 61404
rect 70364 61348 70420 63084
rect 70476 62356 70532 63532
rect 70812 63476 70868 64428
rect 70924 64148 70980 64652
rect 71260 64708 71316 64718
rect 71260 64614 71316 64652
rect 71484 64594 71540 64876
rect 71932 64820 71988 65214
rect 71708 64764 71988 64820
rect 72044 64932 72100 64942
rect 72044 64818 72100 64876
rect 72044 64766 72046 64818
rect 72098 64766 72100 64818
rect 71484 64542 71486 64594
rect 71538 64542 71540 64594
rect 71484 64530 71540 64542
rect 71596 64708 71652 64718
rect 70924 64146 71204 64148
rect 70924 64094 70926 64146
rect 70978 64094 71204 64146
rect 70924 64092 71204 64094
rect 70924 64082 70980 64092
rect 70476 62290 70532 62300
rect 70588 63420 70868 63476
rect 70924 63700 70980 63710
rect 70588 61794 70644 63420
rect 70588 61742 70590 61794
rect 70642 61742 70644 61794
rect 70588 61730 70644 61742
rect 70700 62914 70756 62926
rect 70700 62862 70702 62914
rect 70754 62862 70756 62914
rect 70476 61460 70532 61470
rect 70476 61366 70532 61404
rect 70252 61292 70420 61348
rect 70252 61012 70308 61292
rect 70700 61236 70756 62862
rect 70924 62244 70980 63644
rect 71036 63588 71092 63598
rect 71036 62692 71092 63532
rect 71036 62626 71092 62636
rect 71036 62356 71092 62394
rect 71036 62290 71092 62300
rect 70924 62132 71092 62188
rect 70700 61170 70756 61180
rect 70252 60956 70532 61012
rect 70140 60806 70196 60844
rect 70476 60898 70532 60956
rect 71036 60900 71092 62132
rect 71148 62132 71204 64092
rect 71372 63922 71428 63934
rect 71372 63870 71374 63922
rect 71426 63870 71428 63922
rect 71372 63700 71428 63870
rect 71372 63634 71428 63644
rect 71596 63364 71652 64652
rect 71148 62066 71204 62076
rect 71260 63308 71652 63364
rect 71708 64148 71764 64764
rect 72044 64754 72100 64766
rect 71708 63924 71764 64092
rect 72156 64148 72212 64158
rect 72268 64148 72324 67564
rect 72492 66164 72548 67790
rect 72828 67732 72884 67742
rect 72828 67730 73108 67732
rect 72828 67678 72830 67730
rect 72882 67678 73108 67730
rect 72828 67676 73108 67678
rect 72828 67666 72884 67676
rect 72492 66098 72548 66108
rect 72716 66946 72772 66958
rect 72716 66894 72718 66946
rect 72770 66894 72772 66946
rect 72604 66052 72660 66062
rect 72604 65958 72660 65996
rect 72716 65604 72772 66894
rect 72604 65548 72772 65604
rect 73052 66386 73108 67676
rect 73052 66334 73054 66386
rect 73106 66334 73108 66386
rect 73052 65604 73108 66334
rect 72604 65492 72660 65548
rect 73052 65538 73108 65548
rect 72156 64146 72324 64148
rect 72156 64094 72158 64146
rect 72210 64094 72324 64146
rect 72156 64092 72324 64094
rect 72492 65436 72604 65492
rect 72044 64036 72100 64046
rect 70476 60846 70478 60898
rect 70530 60846 70532 60898
rect 70476 60834 70532 60846
rect 70588 60898 71092 60900
rect 70588 60846 71038 60898
rect 71090 60846 71092 60898
rect 70588 60844 71092 60846
rect 70028 60722 70084 60732
rect 70588 60676 70644 60844
rect 71036 60834 71092 60844
rect 71148 61572 71204 61582
rect 69916 60050 69972 60060
rect 70364 60620 70644 60676
rect 70364 60004 70420 60620
rect 69804 59838 69806 59890
rect 69858 59838 69860 59890
rect 69804 59826 69860 59838
rect 70028 59948 70420 60004
rect 69468 58258 69524 58268
rect 69580 58660 69636 58670
rect 69580 57874 69636 58604
rect 69580 57822 69582 57874
rect 69634 57822 69636 57874
rect 69580 57810 69636 57822
rect 69804 58658 69860 58670
rect 69804 58606 69806 58658
rect 69858 58606 69860 58658
rect 69804 58210 69860 58606
rect 69804 58158 69806 58210
rect 69858 58158 69860 58210
rect 69692 57204 69748 57214
rect 69692 56866 69748 57148
rect 69692 56814 69694 56866
rect 69746 56814 69748 56866
rect 69692 56802 69748 56814
rect 69356 56642 69412 56654
rect 69356 56590 69358 56642
rect 69410 56590 69412 56642
rect 69356 56084 69412 56590
rect 69356 56018 69412 56028
rect 69804 55468 69860 58158
rect 70028 57874 70084 59948
rect 70252 59780 70308 59790
rect 70252 58772 70308 59724
rect 70364 59218 70420 59948
rect 70700 60564 70756 60574
rect 70476 59890 70532 59902
rect 70476 59838 70478 59890
rect 70530 59838 70532 59890
rect 70476 59780 70532 59838
rect 70476 59714 70532 59724
rect 70588 59556 70644 59566
rect 70588 59442 70644 59500
rect 70588 59390 70590 59442
rect 70642 59390 70644 59442
rect 70588 59378 70644 59390
rect 70364 59166 70366 59218
rect 70418 59166 70420 59218
rect 70364 59154 70420 59166
rect 70476 59108 70532 59118
rect 70252 58716 70420 58772
rect 70252 58548 70308 58558
rect 70252 58454 70308 58492
rect 70028 57822 70030 57874
rect 70082 57822 70084 57874
rect 70028 57810 70084 57822
rect 70140 57988 70196 57998
rect 70140 57204 70196 57932
rect 70364 57876 70420 58716
rect 70364 57744 70420 57820
rect 70140 56978 70196 57148
rect 70140 56926 70142 56978
rect 70194 56926 70196 56978
rect 70140 56914 70196 56926
rect 69244 55412 69412 55468
rect 68684 49746 68740 49756
rect 68796 55074 68852 55086
rect 68796 55022 68798 55074
rect 68850 55022 68852 55074
rect 68796 50820 68852 55022
rect 69132 54626 69188 54638
rect 69132 54574 69134 54626
rect 69186 54574 69188 54626
rect 69132 52164 69188 54574
rect 69244 53508 69300 53518
rect 69244 53414 69300 53452
rect 69132 52098 69188 52108
rect 68796 50764 69300 50820
rect 68684 49252 68740 49262
rect 68684 49026 68740 49196
rect 68684 48974 68686 49026
rect 68738 48974 68740 49026
rect 68684 48962 68740 48974
rect 68796 49028 68852 50764
rect 69244 50706 69300 50764
rect 69244 50654 69246 50706
rect 69298 50654 69300 50706
rect 69244 50642 69300 50654
rect 69356 50428 69412 55412
rect 69692 55412 69860 55468
rect 69468 54628 69524 54638
rect 69468 54534 69524 54572
rect 69580 53618 69636 53630
rect 69580 53566 69582 53618
rect 69634 53566 69636 53618
rect 69468 53506 69524 53518
rect 69468 53454 69470 53506
rect 69522 53454 69524 53506
rect 69468 52834 69524 53454
rect 69580 53396 69636 53566
rect 69580 53330 69636 53340
rect 69468 52782 69470 52834
rect 69522 52782 69524 52834
rect 69468 52770 69524 52782
rect 69692 50596 69748 55412
rect 69916 54628 69972 54638
rect 69916 54534 69972 54572
rect 70364 53618 70420 53630
rect 70364 53566 70366 53618
rect 70418 53566 70420 53618
rect 70028 53506 70084 53518
rect 70028 53454 70030 53506
rect 70082 53454 70084 53506
rect 70028 52612 70084 53454
rect 70028 52546 70084 52556
rect 70252 53506 70308 53518
rect 70252 53454 70254 53506
rect 70306 53454 70308 53506
rect 70252 52388 70308 53454
rect 70364 53508 70420 53566
rect 70364 53442 70420 53452
rect 70364 53172 70420 53182
rect 70364 53078 70420 53116
rect 69804 52332 70308 52388
rect 69804 52274 69860 52332
rect 69804 52222 69806 52274
rect 69858 52222 69860 52274
rect 69804 52210 69860 52222
rect 70028 51268 70084 52332
rect 70140 52164 70196 52174
rect 70140 52070 70196 52108
rect 70140 51268 70196 51278
rect 70028 51266 70196 51268
rect 70028 51214 70142 51266
rect 70194 51214 70196 51266
rect 70028 51212 70196 51214
rect 70140 51202 70196 51212
rect 70476 50596 70532 59052
rect 70700 58324 70756 60508
rect 70812 60004 70868 60014
rect 70812 59890 70868 59948
rect 70812 59838 70814 59890
rect 70866 59838 70868 59890
rect 70812 58660 70868 59838
rect 70812 58594 70868 58604
rect 70924 59556 70980 59566
rect 70812 58324 70868 58334
rect 70700 58322 70868 58324
rect 70700 58270 70814 58322
rect 70866 58270 70868 58322
rect 70700 58268 70868 58270
rect 70812 58258 70868 58268
rect 70588 57540 70644 57550
rect 70588 56980 70644 57484
rect 70812 57540 70868 57550
rect 70812 57446 70868 57484
rect 70588 56886 70644 56924
rect 70924 56420 70980 59500
rect 71148 59442 71204 61516
rect 71148 59390 71150 59442
rect 71202 59390 71204 59442
rect 71148 59378 71204 59390
rect 71260 59220 71316 63308
rect 71708 63252 71764 63868
rect 71932 63924 71988 63934
rect 71932 63830 71988 63868
rect 72044 63588 72100 63980
rect 72156 63924 72212 64092
rect 72380 64036 72436 64046
rect 72380 63942 72436 63980
rect 72156 63858 72212 63868
rect 71484 63196 71764 63252
rect 71932 63532 72100 63588
rect 72268 63812 72324 63822
rect 71484 63140 71540 63196
rect 71932 63140 71988 63532
rect 71372 63138 71540 63140
rect 71372 63086 71486 63138
rect 71538 63086 71540 63138
rect 71372 63084 71540 63086
rect 71372 62020 71428 63084
rect 71484 63074 71540 63084
rect 71596 63138 71988 63140
rect 71596 63086 71934 63138
rect 71986 63086 71988 63138
rect 71596 63084 71988 63086
rect 71484 62244 71540 62254
rect 71484 62150 71540 62188
rect 71372 61964 71540 62020
rect 71372 60900 71428 60910
rect 71372 60806 71428 60844
rect 71484 60564 71540 61964
rect 71596 61682 71652 63084
rect 71932 63074 71988 63084
rect 72044 63362 72100 63374
rect 72044 63310 72046 63362
rect 72098 63310 72100 63362
rect 71708 62914 71764 62926
rect 71708 62862 71710 62914
rect 71762 62862 71764 62914
rect 71708 62132 71764 62862
rect 71932 62692 71988 62702
rect 71932 62356 71988 62636
rect 72044 62580 72100 63310
rect 72156 63140 72212 63150
rect 72268 63140 72324 63756
rect 72156 63138 72324 63140
rect 72156 63086 72158 63138
rect 72210 63086 72324 63138
rect 72156 63084 72324 63086
rect 72156 63074 72212 63084
rect 72044 62524 72212 62580
rect 72044 62356 72100 62366
rect 71932 62354 72100 62356
rect 71932 62302 72046 62354
rect 72098 62302 72100 62354
rect 71932 62300 72100 62302
rect 72044 62290 72100 62300
rect 71708 62066 71764 62076
rect 71596 61630 71598 61682
rect 71650 61630 71652 61682
rect 71596 61618 71652 61630
rect 72156 61124 72212 62524
rect 72492 62354 72548 65436
rect 72604 65426 72660 65436
rect 72716 65380 72772 65390
rect 72716 65286 72772 65324
rect 72716 64148 72772 64158
rect 73164 64148 73220 77868
rect 73276 77858 73332 77868
rect 73948 77252 74004 77980
rect 73724 77196 73948 77252
rect 73724 76466 73780 77196
rect 73948 77186 74004 77196
rect 73724 76414 73726 76466
rect 73778 76414 73780 76466
rect 73724 76402 73780 76414
rect 73724 76244 73780 76254
rect 73388 75796 73444 75806
rect 73388 75702 73444 75740
rect 73724 75794 73780 76188
rect 73724 75742 73726 75794
rect 73778 75742 73780 75794
rect 73724 75684 73780 75742
rect 73724 75618 73780 75628
rect 73724 74900 73780 74910
rect 73724 74786 73780 74844
rect 73724 74734 73726 74786
rect 73778 74734 73780 74786
rect 73500 74676 73556 74686
rect 73276 74004 73332 74014
rect 73276 71876 73332 73948
rect 73388 73218 73444 73230
rect 73388 73166 73390 73218
rect 73442 73166 73444 73218
rect 73388 71988 73444 73166
rect 73500 72658 73556 74620
rect 73724 74004 73780 74734
rect 73724 73938 73780 73948
rect 73724 73332 73780 73342
rect 73724 73330 74004 73332
rect 73724 73278 73726 73330
rect 73778 73278 74004 73330
rect 73724 73276 74004 73278
rect 73724 73266 73780 73276
rect 73500 72606 73502 72658
rect 73554 72606 73556 72658
rect 73500 72594 73556 72606
rect 73948 72546 74004 73276
rect 73948 72494 73950 72546
rect 74002 72494 74004 72546
rect 73836 72100 73892 72110
rect 73612 71988 73668 71998
rect 73388 71932 73612 71988
rect 73276 71820 73556 71876
rect 73276 71652 73332 71662
rect 73276 71558 73332 71596
rect 73276 70980 73332 70990
rect 73276 69410 73332 70924
rect 73276 69358 73278 69410
rect 73330 69358 73332 69410
rect 73276 67956 73332 69358
rect 73388 70082 73444 70094
rect 73388 70030 73390 70082
rect 73442 70030 73444 70082
rect 73388 68292 73444 70030
rect 73500 68740 73556 71820
rect 73612 68852 73668 71932
rect 73836 71986 73892 72044
rect 73836 71934 73838 71986
rect 73890 71934 73892 71986
rect 73836 71764 73892 71934
rect 73948 71764 74004 72494
rect 73836 71708 74004 71764
rect 73836 71652 73892 71708
rect 73836 71586 73892 71596
rect 74060 70082 74116 70094
rect 74060 70030 74062 70082
rect 74114 70030 74116 70082
rect 74060 69300 74116 70030
rect 74060 69234 74116 69244
rect 73948 69186 74004 69198
rect 73948 69134 73950 69186
rect 74002 69134 74004 69186
rect 73724 68852 73780 68862
rect 73612 68850 73780 68852
rect 73612 68798 73726 68850
rect 73778 68798 73780 68850
rect 73612 68796 73780 68798
rect 73500 68674 73556 68684
rect 73724 68740 73780 68796
rect 73780 68684 73892 68740
rect 73724 68674 73780 68684
rect 73388 68226 73444 68236
rect 73724 68292 73780 68302
rect 73388 67956 73444 67966
rect 73276 67954 73444 67956
rect 73276 67902 73390 67954
rect 73442 67902 73444 67954
rect 73276 67900 73444 67902
rect 73388 67890 73444 67900
rect 73388 67396 73444 67406
rect 73388 67282 73444 67340
rect 73388 67230 73390 67282
rect 73442 67230 73444 67282
rect 73388 67218 73444 67230
rect 73500 66948 73556 66958
rect 72716 64146 73220 64148
rect 72716 64094 72718 64146
rect 72770 64094 73220 64146
rect 72716 64092 73220 64094
rect 73276 66052 73332 66062
rect 73276 64594 73332 65996
rect 73500 65714 73556 66892
rect 73724 66836 73780 68236
rect 73836 67844 73892 68684
rect 73948 68180 74004 69134
rect 73948 68114 74004 68124
rect 74060 69076 74116 69086
rect 73836 67712 73892 67788
rect 73948 67172 74004 67182
rect 73948 66948 74004 67116
rect 73612 66834 73780 66836
rect 73612 66782 73726 66834
rect 73778 66782 73780 66834
rect 73612 66780 73780 66782
rect 73612 66052 73668 66780
rect 73724 66770 73780 66780
rect 73836 66892 74004 66948
rect 73724 66164 73780 66174
rect 73836 66164 73892 66892
rect 74060 66498 74116 69020
rect 74060 66446 74062 66498
rect 74114 66446 74116 66498
rect 74060 66434 74116 66446
rect 74060 66276 74116 66286
rect 74060 66182 74116 66220
rect 73780 66108 73892 66164
rect 73724 66070 73780 66108
rect 73612 65986 73668 65996
rect 73500 65662 73502 65714
rect 73554 65662 73556 65714
rect 73500 65650 73556 65662
rect 73948 65602 74004 65614
rect 73948 65550 73950 65602
rect 74002 65550 74004 65602
rect 73948 65492 74004 65550
rect 73276 64542 73278 64594
rect 73330 64542 73332 64594
rect 72716 64082 72772 64092
rect 72604 63922 72660 63934
rect 72604 63870 72606 63922
rect 72658 63870 72660 63922
rect 72604 63812 72660 63870
rect 72604 63746 72660 63756
rect 72716 63924 72772 63934
rect 72492 62302 72494 62354
rect 72546 62302 72548 62354
rect 72492 62188 72548 62302
rect 72716 63138 72772 63868
rect 72716 63086 72718 63138
rect 72770 63086 72772 63138
rect 72716 62188 72772 63086
rect 72380 62132 72548 62188
rect 72604 62132 72772 62188
rect 72380 61908 72436 62132
rect 72380 61842 72436 61852
rect 72492 62020 72548 62030
rect 72492 61684 72548 61964
rect 72380 61682 72548 61684
rect 72380 61630 72494 61682
rect 72546 61630 72548 61682
rect 72380 61628 72548 61630
rect 71484 60498 71540 60508
rect 72044 61068 72212 61124
rect 72268 61572 72324 61582
rect 71484 60114 71540 60126
rect 71484 60062 71486 60114
rect 71538 60062 71540 60114
rect 71484 59332 71540 60062
rect 71932 60004 71988 60014
rect 71932 59910 71988 59948
rect 72044 59444 72100 61068
rect 72156 60900 72212 60910
rect 72156 60786 72212 60844
rect 72156 60734 72158 60786
rect 72210 60734 72212 60786
rect 72156 60722 72212 60734
rect 70924 56306 70980 56364
rect 70924 56254 70926 56306
rect 70978 56254 70980 56306
rect 70924 56242 70980 56254
rect 71036 59164 71316 59220
rect 71372 59218 71428 59230
rect 71372 59166 71374 59218
rect 71426 59166 71428 59218
rect 70700 55298 70756 55310
rect 70700 55246 70702 55298
rect 70754 55246 70756 55298
rect 70700 54628 70756 55246
rect 70700 54562 70756 54572
rect 70924 55074 70980 55086
rect 70924 55022 70926 55074
rect 70978 55022 70980 55074
rect 70812 53506 70868 53518
rect 70812 53454 70814 53506
rect 70866 53454 70868 53506
rect 70812 53396 70868 53454
rect 70924 53508 70980 55022
rect 70924 53442 70980 53452
rect 70812 53330 70868 53340
rect 70812 53058 70868 53070
rect 70812 53006 70814 53058
rect 70866 53006 70868 53058
rect 70812 52388 70868 53006
rect 70812 52322 70868 52332
rect 70700 52162 70756 52174
rect 70700 52110 70702 52162
rect 70754 52110 70756 52162
rect 70700 52052 70756 52110
rect 70700 51986 70756 51996
rect 70812 52052 70868 52062
rect 71036 52052 71092 59164
rect 71372 58772 71428 59166
rect 71148 58322 71204 58334
rect 71148 58270 71150 58322
rect 71202 58270 71204 58322
rect 71148 57092 71204 58270
rect 71372 57540 71428 58716
rect 71484 58660 71540 59276
rect 71484 58594 71540 58604
rect 71932 59388 72100 59444
rect 72156 60564 72212 60574
rect 71596 58324 71652 58334
rect 71596 57652 71652 58268
rect 71820 58324 71876 58362
rect 71820 58258 71876 58268
rect 71932 58212 71988 59388
rect 72044 59218 72100 59230
rect 72044 59166 72046 59218
rect 72098 59166 72100 59218
rect 72044 58772 72100 59166
rect 72156 58828 72212 60508
rect 72268 60340 72324 61516
rect 72268 60274 72324 60284
rect 72156 58772 72324 58828
rect 72044 58706 72100 58716
rect 72268 58546 72324 58772
rect 72268 58494 72270 58546
rect 72322 58494 72324 58546
rect 72268 58482 72324 58494
rect 72156 58434 72212 58446
rect 72156 58382 72158 58434
rect 72210 58382 72212 58434
rect 72156 58212 72212 58382
rect 71932 58156 72100 58212
rect 71820 58100 71876 58110
rect 71596 57650 71764 57652
rect 71596 57598 71598 57650
rect 71650 57598 71764 57650
rect 71596 57596 71764 57598
rect 71596 57586 71652 57596
rect 71372 57474 71428 57484
rect 71148 57026 71204 57036
rect 71708 56868 71764 57596
rect 71820 57650 71876 58044
rect 71820 57598 71822 57650
rect 71874 57598 71876 57650
rect 71820 57586 71876 57598
rect 71820 56868 71876 56878
rect 71708 56866 71876 56868
rect 71708 56814 71822 56866
rect 71874 56814 71876 56866
rect 71708 56812 71876 56814
rect 71820 56802 71876 56812
rect 71148 56644 71204 56654
rect 71148 56550 71204 56588
rect 71596 56642 71652 56654
rect 71596 56590 71598 56642
rect 71650 56590 71652 56642
rect 71484 56532 71540 56542
rect 71484 56306 71540 56476
rect 71484 56254 71486 56306
rect 71538 56254 71540 56306
rect 71484 56242 71540 56254
rect 71596 55468 71652 56590
rect 72044 56532 72100 58156
rect 72156 58146 72212 58156
rect 71932 56308 71988 56318
rect 71932 56214 71988 56252
rect 71596 55412 71764 55468
rect 71148 54628 71204 54638
rect 71148 54534 71204 54572
rect 71708 54402 71764 55412
rect 72044 55298 72100 56476
rect 72156 57426 72212 57438
rect 72156 57374 72158 57426
rect 72210 57374 72212 57426
rect 72156 57092 72212 57374
rect 72380 57092 72436 61628
rect 72492 61618 72548 61628
rect 72492 60900 72548 60910
rect 72492 60002 72548 60844
rect 72604 60900 72660 62132
rect 72828 61908 72884 61918
rect 72828 61460 72884 61852
rect 72828 61366 72884 61404
rect 73276 61908 73332 64542
rect 72940 61236 72996 61246
rect 72604 60898 72884 60900
rect 72604 60846 72606 60898
rect 72658 60846 72884 60898
rect 72604 60844 72884 60846
rect 72604 60834 72660 60844
rect 72716 60340 72772 60350
rect 72716 60226 72772 60284
rect 72716 60174 72718 60226
rect 72770 60174 72772 60226
rect 72716 60162 72772 60174
rect 72492 59950 72494 60002
rect 72546 59950 72548 60002
rect 72492 59938 72548 59950
rect 72604 60004 72660 60014
rect 72604 59218 72660 59948
rect 72604 59166 72606 59218
rect 72658 59166 72660 59218
rect 72604 59154 72660 59166
rect 72828 58436 72884 60844
rect 72940 60228 72996 61180
rect 73276 60564 73332 61852
rect 73724 65380 73780 65390
rect 73724 61572 73780 65324
rect 73948 64036 74004 65436
rect 73836 64034 74004 64036
rect 73836 63982 73950 64034
rect 74002 63982 74004 64034
rect 73836 63980 74004 63982
rect 73836 63026 73892 63980
rect 73948 63904 74004 63980
rect 74060 64708 74116 64718
rect 73836 62974 73838 63026
rect 73890 62974 73892 63026
rect 73836 62962 73892 62974
rect 74060 62244 74116 64652
rect 74172 64482 74228 78652
rect 74620 77924 74676 77934
rect 74620 77922 74788 77924
rect 74620 77870 74622 77922
rect 74674 77870 74788 77922
rect 74620 77868 74788 77870
rect 74620 77858 74676 77868
rect 74732 77140 74788 77868
rect 74956 77812 75012 80220
rect 74956 77746 75012 77756
rect 74732 77074 74788 77084
rect 74956 77138 75012 77150
rect 74956 77086 74958 77138
rect 75010 77086 75012 77138
rect 74284 77028 74340 77038
rect 74620 77028 74676 77038
rect 74284 76244 74340 76972
rect 74396 77026 74676 77028
rect 74396 76974 74622 77026
rect 74674 76974 74676 77026
rect 74396 76972 74676 76974
rect 74396 76578 74452 76972
rect 74620 76962 74676 76972
rect 74844 77026 74900 77038
rect 74844 76974 74846 77026
rect 74898 76974 74900 77026
rect 74396 76526 74398 76578
rect 74450 76526 74452 76578
rect 74396 76514 74452 76526
rect 74284 76178 74340 76188
rect 74396 76356 74452 76366
rect 74284 75796 74340 75806
rect 74284 75570 74340 75740
rect 74284 75518 74286 75570
rect 74338 75518 74340 75570
rect 74284 75506 74340 75518
rect 74396 75458 74452 76300
rect 74844 76020 74900 76974
rect 74620 75964 74900 76020
rect 74620 75682 74676 75964
rect 74620 75630 74622 75682
rect 74674 75630 74676 75682
rect 74620 75618 74676 75630
rect 74956 75684 75012 77086
rect 75068 75796 75124 81116
rect 75180 80500 75236 80510
rect 75180 80274 75236 80444
rect 75292 80386 75348 81340
rect 75292 80334 75294 80386
rect 75346 80334 75348 80386
rect 75292 80322 75348 80334
rect 75180 80222 75182 80274
rect 75234 80222 75236 80274
rect 75180 80210 75236 80222
rect 75404 78988 75460 81564
rect 75964 80612 76020 80622
rect 75292 78932 75460 78988
rect 75740 80162 75796 80174
rect 75740 80110 75742 80162
rect 75794 80110 75796 80162
rect 75180 78708 75236 78718
rect 75180 78614 75236 78652
rect 75068 75740 75236 75796
rect 74956 75618 75012 75628
rect 75068 75572 75124 75582
rect 75068 75478 75124 75516
rect 74396 75406 74398 75458
rect 74450 75406 74452 75458
rect 74396 75012 74452 75406
rect 74620 75124 74676 75134
rect 74620 75030 74676 75068
rect 74396 74946 74452 74956
rect 75068 75012 75124 75022
rect 75068 74918 75124 74956
rect 74284 74900 74340 74910
rect 74284 74806 74340 74844
rect 75180 74340 75236 75740
rect 74732 74284 75236 74340
rect 74396 73330 74452 73342
rect 74396 73278 74398 73330
rect 74450 73278 74452 73330
rect 74396 72212 74452 73278
rect 74396 72146 74452 72156
rect 74284 71650 74340 71662
rect 74284 71598 74286 71650
rect 74338 71598 74340 71650
rect 74284 71204 74340 71598
rect 74284 71138 74340 71148
rect 74732 69076 74788 74284
rect 74844 74114 74900 74126
rect 74844 74062 74846 74114
rect 74898 74062 74900 74114
rect 74844 72770 74900 74062
rect 75068 73890 75124 73902
rect 75068 73838 75070 73890
rect 75122 73838 75124 73890
rect 75068 73442 75124 73838
rect 75068 73390 75070 73442
rect 75122 73390 75124 73442
rect 75068 73378 75124 73390
rect 74844 72718 74846 72770
rect 74898 72718 74900 72770
rect 74844 72706 74900 72718
rect 75180 72548 75236 72558
rect 75292 72548 75348 78932
rect 75740 78820 75796 80110
rect 75740 78754 75796 78764
rect 75964 78818 76020 80556
rect 76188 80164 76244 80174
rect 76188 80070 76244 80108
rect 77196 79716 77252 81676
rect 77308 81666 77364 81676
rect 78316 80724 78372 82574
rect 78316 80658 78372 80668
rect 77196 79660 77364 79716
rect 76300 79492 76356 79502
rect 75964 78766 75966 78818
rect 76018 78766 76020 78818
rect 75964 78754 76020 78766
rect 76188 79490 76356 79492
rect 76188 79438 76302 79490
rect 76354 79438 76356 79490
rect 76188 79436 76356 79438
rect 75516 78708 75572 78718
rect 75516 78614 75572 78652
rect 76188 78594 76244 79436
rect 76300 79426 76356 79436
rect 76748 79490 76804 79502
rect 77196 79492 77252 79502
rect 76748 79438 76750 79490
rect 76802 79438 76804 79490
rect 76300 78708 76356 78718
rect 76300 78614 76356 78652
rect 76748 78708 76804 79438
rect 76748 78642 76804 78652
rect 76972 79436 77196 79492
rect 76188 78542 76190 78594
rect 76242 78542 76244 78594
rect 76188 78148 76244 78542
rect 76188 78082 76244 78092
rect 76748 78036 76804 78046
rect 76748 77922 76804 77980
rect 76748 77870 76750 77922
rect 76802 77870 76804 77922
rect 76748 77858 76804 77870
rect 76524 77252 76580 77262
rect 76524 77158 76580 77196
rect 76972 77252 77028 79436
rect 77196 79398 77252 79436
rect 77308 79268 77364 79660
rect 75516 77138 75572 77150
rect 75516 77086 75518 77138
rect 75570 77086 75572 77138
rect 75516 77028 75572 77086
rect 75516 76962 75572 76972
rect 75852 77026 75908 77038
rect 75852 76974 75854 77026
rect 75906 76974 75908 77026
rect 75852 76692 75908 76974
rect 75852 76626 75908 76636
rect 76972 76690 77028 77196
rect 76972 76638 76974 76690
rect 77026 76638 77028 76690
rect 76972 76626 77028 76638
rect 77084 79212 77364 79268
rect 75404 76580 75460 76590
rect 75404 75796 75460 76524
rect 76524 76356 76580 76366
rect 75404 75570 75460 75740
rect 76076 76354 76580 76356
rect 76076 76302 76526 76354
rect 76578 76302 76580 76354
rect 76076 76300 76580 76302
rect 75404 75518 75406 75570
rect 75458 75518 75460 75570
rect 75404 75506 75460 75518
rect 75964 75572 76020 75582
rect 75964 75124 76020 75516
rect 76076 75570 76132 76300
rect 76524 76290 76580 76300
rect 76300 75684 76356 75694
rect 76300 75590 76356 75628
rect 76076 75518 76078 75570
rect 76130 75518 76132 75570
rect 76076 75506 76132 75518
rect 76076 75124 76132 75134
rect 76020 75122 76132 75124
rect 76020 75070 76078 75122
rect 76130 75070 76132 75122
rect 76020 75068 76132 75070
rect 75964 74992 76020 75068
rect 76076 75058 76132 75068
rect 75740 74786 75796 74798
rect 75740 74734 75742 74786
rect 75794 74734 75796 74786
rect 75740 74116 75796 74734
rect 76076 74116 76132 74126
rect 75740 74114 76132 74116
rect 75740 74062 76078 74114
rect 76130 74062 76132 74114
rect 75740 74060 76132 74062
rect 75964 73220 76020 73230
rect 75180 72546 75348 72548
rect 75180 72494 75182 72546
rect 75234 72494 75348 72546
rect 75180 72492 75348 72494
rect 75628 72546 75684 72558
rect 75628 72494 75630 72546
rect 75682 72494 75684 72546
rect 75180 72324 75236 72492
rect 75180 72258 75236 72268
rect 75628 72100 75684 72494
rect 75964 72434 76020 73164
rect 75964 72382 75966 72434
rect 76018 72382 76020 72434
rect 75964 72370 76020 72382
rect 74844 71988 74900 71998
rect 74844 71650 74900 71932
rect 74844 71598 74846 71650
rect 74898 71598 74900 71650
rect 74844 71538 74900 71598
rect 74844 71486 74846 71538
rect 74898 71486 74900 71538
rect 74844 71474 74900 71486
rect 75068 71652 75124 71662
rect 74956 69412 75012 69422
rect 74844 69300 74900 69310
rect 74844 69206 74900 69244
rect 74732 69010 74788 69020
rect 74284 68852 74340 68862
rect 74284 68628 74340 68796
rect 74844 68852 74900 68862
rect 74956 68852 75012 69356
rect 74844 68850 75012 68852
rect 74844 68798 74846 68850
rect 74898 68798 75012 68850
rect 74844 68796 75012 68798
rect 74844 68786 74900 68796
rect 74284 68496 74340 68572
rect 74844 68404 74900 68414
rect 75068 68404 75124 71596
rect 75292 71650 75348 71662
rect 75292 71598 75294 71650
rect 75346 71598 75348 71650
rect 75292 71538 75348 71598
rect 75292 71486 75294 71538
rect 75346 71486 75348 71538
rect 75292 71474 75348 71486
rect 75628 71204 75684 72044
rect 75628 71138 75684 71148
rect 75740 71650 75796 71662
rect 75740 71598 75742 71650
rect 75794 71598 75796 71650
rect 75292 70978 75348 70990
rect 75292 70926 75294 70978
rect 75346 70926 75348 70978
rect 75180 69860 75236 69870
rect 75180 69298 75236 69804
rect 75292 69636 75348 70926
rect 75516 70754 75572 70766
rect 75516 70702 75518 70754
rect 75570 70702 75572 70754
rect 75516 70308 75572 70702
rect 75516 70242 75572 70252
rect 75740 69860 75796 71598
rect 76076 71652 76132 74060
rect 76524 74114 76580 74126
rect 76524 74062 76526 74114
rect 76578 74062 76580 74114
rect 76524 73444 76580 74062
rect 77084 73948 77140 79212
rect 78428 78988 78484 90692
rect 81276 89404 81540 89414
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81276 89338 81540 89348
rect 81276 87836 81540 87846
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81276 87770 81540 87780
rect 81788 86884 81844 86894
rect 81788 86882 82068 86884
rect 81788 86830 81790 86882
rect 81842 86830 82068 86882
rect 81788 86828 82068 86830
rect 81788 86818 81844 86828
rect 81900 86546 81956 86558
rect 81900 86494 81902 86546
rect 81954 86494 81956 86546
rect 78652 86434 78708 86446
rect 78652 86382 78654 86434
rect 78706 86382 78708 86434
rect 78652 85986 78708 86382
rect 79660 86434 79716 86446
rect 79660 86382 79662 86434
rect 79714 86382 79716 86434
rect 79212 86100 79268 86110
rect 79212 86006 79268 86044
rect 78652 85934 78654 85986
rect 78706 85934 78708 85986
rect 78540 83412 78596 83422
rect 78540 83318 78596 83356
rect 78652 82068 78708 85934
rect 78876 85764 78932 85774
rect 78876 85670 78932 85708
rect 79660 85764 79716 86382
rect 81228 86436 81284 86474
rect 81788 86436 81844 86446
rect 81228 86370 81284 86380
rect 81676 86434 81844 86436
rect 81676 86382 81790 86434
rect 81842 86382 81844 86434
rect 81676 86380 81844 86382
rect 81276 86268 81540 86278
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81276 86202 81540 86212
rect 81676 86100 81732 86380
rect 81788 86370 81844 86380
rect 81900 86436 81956 86494
rect 81900 86370 81956 86380
rect 81340 86044 81732 86100
rect 78764 84978 78820 84990
rect 78764 84926 78766 84978
rect 78818 84926 78820 84978
rect 78764 84308 78820 84926
rect 78764 82962 78820 84252
rect 79548 84308 79604 84318
rect 79548 83634 79604 84252
rect 79660 84196 79716 85708
rect 79772 85762 79828 85774
rect 79772 85710 79774 85762
rect 79826 85710 79828 85762
rect 79772 85652 79828 85710
rect 79772 85586 79828 85596
rect 80444 85762 80500 85774
rect 80444 85710 80446 85762
rect 80498 85710 80500 85762
rect 80444 85652 80500 85710
rect 81340 85762 81396 86044
rect 81340 85710 81342 85762
rect 81394 85710 81396 85762
rect 81340 85698 81396 85710
rect 80444 84308 80500 85596
rect 81676 85652 81732 85662
rect 81276 84700 81540 84710
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81276 84634 81540 84644
rect 81676 84420 81732 85596
rect 80332 84252 80444 84308
rect 80220 84196 80276 84206
rect 79660 84194 80276 84196
rect 79660 84142 80222 84194
rect 80274 84142 80276 84194
rect 79660 84140 80276 84142
rect 79548 83582 79550 83634
rect 79602 83582 79604 83634
rect 79548 83570 79604 83582
rect 78764 82910 78766 82962
rect 78818 82910 78820 82962
rect 78764 82898 78820 82910
rect 79212 83298 79268 83310
rect 79212 83246 79214 83298
rect 79266 83246 79268 83298
rect 79212 82292 79268 83246
rect 80108 83300 80164 84140
rect 80220 84130 80276 84140
rect 80220 83524 80276 83534
rect 80332 83524 80388 84252
rect 80444 84242 80500 84252
rect 81452 84308 81508 84318
rect 81452 84214 81508 84252
rect 80220 83522 80388 83524
rect 80220 83470 80222 83522
rect 80274 83470 80388 83522
rect 80220 83468 80388 83470
rect 80556 84196 80612 84206
rect 80220 83458 80276 83468
rect 80444 83412 80500 83422
rect 80108 83244 80276 83300
rect 79212 82226 79268 82236
rect 78652 82002 78708 82012
rect 80108 81172 80164 81182
rect 80108 81078 80164 81116
rect 79548 80948 79604 80958
rect 79324 80724 79380 80734
rect 78876 80386 78932 80398
rect 78876 80334 78878 80386
rect 78930 80334 78932 80386
rect 78876 79492 78932 80334
rect 78876 79044 78932 79436
rect 78932 78988 79044 79044
rect 78428 78932 78708 78988
rect 78876 78978 78932 78988
rect 77308 78148 77364 78158
rect 77308 78054 77364 78092
rect 78316 78148 78372 78158
rect 78316 78146 78484 78148
rect 78316 78094 78318 78146
rect 78370 78094 78484 78146
rect 78316 78092 78484 78094
rect 78316 78082 78372 78092
rect 77756 78034 77812 78046
rect 77756 77982 77758 78034
rect 77810 77982 77812 78034
rect 77756 77364 77812 77982
rect 77756 77298 77812 77308
rect 78092 78036 78148 78046
rect 77196 77140 77252 77150
rect 77196 77046 77252 77084
rect 77532 77140 77588 77150
rect 77980 77140 78036 77150
rect 77532 77138 78036 77140
rect 77532 77086 77534 77138
rect 77586 77086 77982 77138
rect 78034 77086 78036 77138
rect 77532 77084 78036 77086
rect 78092 77140 78148 77980
rect 78316 77252 78372 77262
rect 78204 77140 78260 77150
rect 78092 77138 78260 77140
rect 78092 77086 78206 77138
rect 78258 77086 78260 77138
rect 78092 77084 78260 77086
rect 77532 77074 77588 77084
rect 77980 77074 78036 77084
rect 78204 77074 78260 77084
rect 78316 77138 78372 77196
rect 78316 77086 78318 77138
rect 78370 77086 78372 77138
rect 77420 77026 77476 77038
rect 77420 76974 77422 77026
rect 77474 76974 77476 77026
rect 77420 75684 77476 76974
rect 77756 76692 77812 76702
rect 77756 76598 77812 76636
rect 78316 76692 78372 77086
rect 78316 76626 78372 76636
rect 77420 75618 77476 75628
rect 78428 74900 78484 78092
rect 78540 77476 78596 77486
rect 78540 76690 78596 77420
rect 78540 76638 78542 76690
rect 78594 76638 78596 76690
rect 78540 76626 78596 76638
rect 78428 74834 78484 74844
rect 76524 73378 76580 73388
rect 76636 73892 77140 73948
rect 77420 74002 77476 74014
rect 77420 73950 77422 74002
rect 77474 73950 77476 74002
rect 76524 72322 76580 72334
rect 76524 72270 76526 72322
rect 76578 72270 76580 72322
rect 76524 72100 76580 72270
rect 76524 72034 76580 72044
rect 76636 71876 76692 73892
rect 77196 73220 77252 73230
rect 77196 73126 77252 73164
rect 77196 72324 77252 72334
rect 77196 72230 77252 72268
rect 77420 72212 77476 73950
rect 78540 74002 78596 74014
rect 78540 73950 78542 74002
rect 78594 73950 78596 74002
rect 78204 73892 78260 73902
rect 78204 73890 78484 73892
rect 78204 73838 78206 73890
rect 78258 73838 78484 73890
rect 78204 73836 78484 73838
rect 78204 73826 78260 73836
rect 77868 73444 77924 73454
rect 77868 72658 77924 73388
rect 78316 73442 78372 73454
rect 78316 73390 78318 73442
rect 78370 73390 78372 73442
rect 78316 73220 78372 73390
rect 78316 73154 78372 73164
rect 77868 72606 77870 72658
rect 77922 72606 77924 72658
rect 77868 72594 77924 72606
rect 77476 72156 77700 72212
rect 77420 72146 77476 72156
rect 76524 71820 76692 71876
rect 76076 71586 76132 71596
rect 76300 71650 76356 71662
rect 76300 71598 76302 71650
rect 76354 71598 76356 71650
rect 76076 70980 76132 70990
rect 76076 70886 76132 70924
rect 76188 70308 76244 70318
rect 76188 70214 76244 70252
rect 75740 69794 75796 69804
rect 75740 69636 75796 69646
rect 75292 69634 75796 69636
rect 75292 69582 75742 69634
rect 75794 69582 75796 69634
rect 75292 69580 75796 69582
rect 75740 69570 75796 69580
rect 76300 69524 76356 71598
rect 76300 69458 76356 69468
rect 76412 70754 76468 70766
rect 76412 70702 76414 70754
rect 76466 70702 76468 70754
rect 75404 69412 75460 69422
rect 75404 69318 75460 69356
rect 75180 69246 75182 69298
rect 75234 69246 75236 69298
rect 75180 68852 75236 69246
rect 76300 69188 76356 69198
rect 75180 68786 75236 68796
rect 76188 69186 76356 69188
rect 76188 69134 76302 69186
rect 76354 69134 76356 69186
rect 76188 69132 76356 69134
rect 75740 68740 75796 68750
rect 75740 68646 75796 68684
rect 75180 68628 75236 68638
rect 75180 68626 75348 68628
rect 75180 68574 75182 68626
rect 75234 68574 75348 68626
rect 75180 68572 75348 68574
rect 75180 68562 75236 68572
rect 75068 68348 75236 68404
rect 74172 64430 74174 64482
rect 74226 64430 74228 64482
rect 74172 64418 74228 64430
rect 74284 67732 74340 67742
rect 74284 64260 74340 67676
rect 74508 67618 74564 67630
rect 74508 67566 74510 67618
rect 74562 67566 74564 67618
rect 74508 67508 74564 67566
rect 74508 67442 74564 67452
rect 74508 67284 74564 67294
rect 74844 67284 74900 68348
rect 74956 67620 75012 67630
rect 75068 67620 75124 67630
rect 74956 67618 75068 67620
rect 74956 67566 74958 67618
rect 75010 67566 75068 67618
rect 74956 67564 75068 67566
rect 74956 67554 75012 67564
rect 74844 67228 75012 67284
rect 74508 67190 74564 67228
rect 74732 67058 74788 67070
rect 74732 67006 74734 67058
rect 74786 67006 74788 67058
rect 74732 66948 74788 67006
rect 74732 66882 74788 66892
rect 74956 66388 75012 67228
rect 74620 66332 75012 66388
rect 74620 66162 74676 66332
rect 74620 66110 74622 66162
rect 74674 66110 74676 66162
rect 74620 66098 74676 66110
rect 74732 66164 74788 66174
rect 74396 64708 74452 64718
rect 74396 64614 74452 64652
rect 73948 61572 74004 61582
rect 73724 61570 74004 61572
rect 73724 61518 73950 61570
rect 74002 61518 74004 61570
rect 73724 61516 74004 61518
rect 73276 60498 73332 60508
rect 73500 60788 73556 60798
rect 72940 60134 72996 60172
rect 73052 59892 73108 59902
rect 73052 59890 73444 59892
rect 73052 59838 73054 59890
rect 73106 59838 73444 59890
rect 73052 59836 73444 59838
rect 73052 59826 73108 59836
rect 72828 58380 72996 58436
rect 72828 58212 72884 58222
rect 72828 58118 72884 58156
rect 72156 56196 72212 57036
rect 72156 56130 72212 56140
rect 72268 57036 72436 57092
rect 72492 57652 72548 57662
rect 72044 55246 72046 55298
rect 72098 55246 72100 55298
rect 72044 55234 72100 55246
rect 71708 54350 71710 54402
rect 71762 54350 71764 54402
rect 71148 53620 71204 53630
rect 71148 53172 71204 53564
rect 71708 53620 71764 54350
rect 71708 53554 71764 53564
rect 71820 55074 71876 55086
rect 71820 55022 71822 55074
rect 71874 55022 71876 55074
rect 71260 53508 71316 53518
rect 71260 53414 71316 53452
rect 71820 53396 71876 55022
rect 72268 54740 72324 57036
rect 72492 56306 72548 57596
rect 72604 57540 72660 57550
rect 72660 57484 72772 57540
rect 72604 57446 72660 57484
rect 72716 56978 72772 57484
rect 72716 56926 72718 56978
rect 72770 56926 72772 56978
rect 72716 56914 72772 56926
rect 72492 56254 72494 56306
rect 72546 56254 72548 56306
rect 72492 56242 72548 56254
rect 72604 56420 72660 56430
rect 72380 56196 72436 56206
rect 72380 56102 72436 56140
rect 72268 54646 72324 54684
rect 72492 55858 72548 55870
rect 72492 55806 72494 55858
rect 72546 55806 72548 55858
rect 72492 53732 72548 55806
rect 72604 54738 72660 56364
rect 72716 56308 72772 56318
rect 72716 55298 72772 56252
rect 72940 56308 72996 58380
rect 73052 58324 73108 58334
rect 73052 56978 73108 58268
rect 73276 58322 73332 58334
rect 73276 58270 73278 58322
rect 73330 58270 73332 58322
rect 73052 56926 73054 56978
rect 73106 56926 73108 56978
rect 73052 56914 73108 56926
rect 73164 57876 73220 57886
rect 72940 56242 72996 56252
rect 73164 55468 73220 57820
rect 72716 55246 72718 55298
rect 72770 55246 72772 55298
rect 72716 55234 72772 55246
rect 73052 55412 73220 55468
rect 72604 54686 72606 54738
rect 72658 54686 72660 54738
rect 72604 53954 72660 54686
rect 72604 53902 72606 53954
rect 72658 53902 72660 53954
rect 72604 53890 72660 53902
rect 72492 53676 72660 53732
rect 71820 53330 71876 53340
rect 72492 53506 72548 53518
rect 72492 53454 72494 53506
rect 72546 53454 72548 53506
rect 71148 53040 71204 53116
rect 72268 53172 72324 53182
rect 72492 53172 72548 53454
rect 72604 53396 72660 53676
rect 73052 53506 73108 55412
rect 73052 53454 73054 53506
rect 73106 53454 73108 53506
rect 72604 53340 72996 53396
rect 72268 53170 72548 53172
rect 72268 53118 72270 53170
rect 72322 53118 72548 53170
rect 72268 53116 72548 53118
rect 72268 53106 72324 53116
rect 72492 52948 72548 53116
rect 72492 52882 72548 52892
rect 71708 52834 71764 52846
rect 71708 52782 71710 52834
rect 71762 52782 71764 52834
rect 71260 52388 71316 52398
rect 71260 52162 71316 52332
rect 71708 52276 71764 52782
rect 71708 52210 71764 52220
rect 72828 52836 72884 52846
rect 71260 52110 71262 52162
rect 71314 52110 71316 52162
rect 71260 52098 71316 52110
rect 72044 52162 72100 52174
rect 72828 52164 72884 52780
rect 72044 52110 72046 52162
rect 72098 52110 72100 52162
rect 70812 52050 71092 52052
rect 70812 51998 70814 52050
rect 70866 51998 71092 52050
rect 70812 51996 71092 51998
rect 70812 51986 70868 51996
rect 72044 51492 72100 52110
rect 72044 51426 72100 51436
rect 72604 52162 72884 52164
rect 72604 52110 72830 52162
rect 72882 52110 72884 52162
rect 72604 52108 72884 52110
rect 72268 51380 72324 51390
rect 69692 50540 69860 50596
rect 69244 50372 69412 50428
rect 69692 50372 69748 50382
rect 68908 49924 68964 49934
rect 68908 49830 68964 49868
rect 68796 48962 68852 48972
rect 68684 48244 68740 48254
rect 68236 48242 68516 48244
rect 68236 48190 68238 48242
rect 68290 48190 68516 48242
rect 68236 48188 68516 48190
rect 68572 48242 68740 48244
rect 68572 48190 68686 48242
rect 68738 48190 68740 48242
rect 68572 48188 68740 48190
rect 68236 48178 68292 48188
rect 67788 47572 67844 47582
rect 67900 47572 67956 47964
rect 67788 47570 67956 47572
rect 67788 47518 67790 47570
rect 67842 47518 67956 47570
rect 67788 47516 67956 47518
rect 67788 47506 67844 47516
rect 68348 47348 68404 47358
rect 67452 46844 67732 46900
rect 68236 47234 68292 47246
rect 68236 47182 68238 47234
rect 68290 47182 68292 47234
rect 67452 46340 67508 46844
rect 67564 46564 67620 46574
rect 67564 46562 68180 46564
rect 67564 46510 67566 46562
rect 67618 46510 68180 46562
rect 67564 46508 68180 46510
rect 67564 46498 67620 46508
rect 67452 46284 67620 46340
rect 67228 44270 67230 44322
rect 67282 44270 67284 44322
rect 67228 44212 67284 44270
rect 67228 42868 67284 44156
rect 67228 42802 67284 42812
rect 67452 45108 67508 45118
rect 66332 41918 66334 41970
rect 66386 41918 66388 41970
rect 66332 41906 66388 41918
rect 66444 42530 66500 42542
rect 66444 42478 66446 42530
rect 66498 42478 66500 42530
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65436 41458 65492 41468
rect 65548 41300 65604 41310
rect 65604 41244 65716 41300
rect 65548 41206 65604 41244
rect 65212 40402 65380 40404
rect 65212 40350 65326 40402
rect 65378 40350 65380 40402
rect 65212 40348 65380 40350
rect 64764 38612 65044 38668
rect 64988 38276 65044 38612
rect 63420 37438 63422 37490
rect 63474 37438 63476 37490
rect 63420 37426 63476 37438
rect 64316 38220 65044 38276
rect 64316 37378 64372 38220
rect 64540 38052 64596 38062
rect 64316 37326 64318 37378
rect 64370 37326 64372 37378
rect 64316 37314 64372 37326
rect 64428 37380 64484 37390
rect 64428 37266 64484 37324
rect 64428 37214 64430 37266
rect 64482 37214 64484 37266
rect 64428 37202 64484 37214
rect 63756 37042 63812 37054
rect 63756 36990 63758 37042
rect 63810 36990 63812 37042
rect 63756 36036 63812 36990
rect 63756 35970 63812 35980
rect 64316 36036 64372 36046
rect 63308 34290 63364 34300
rect 63644 35586 63700 35598
rect 63644 35534 63646 35586
rect 63698 35534 63700 35586
rect 63644 35028 63700 35534
rect 62076 33628 62244 33684
rect 62076 33458 62132 33628
rect 62076 33406 62078 33458
rect 62130 33406 62132 33458
rect 62076 33394 62132 33406
rect 63532 32788 63588 32798
rect 63644 32788 63700 34972
rect 64316 35026 64372 35980
rect 64540 35922 64596 37996
rect 64876 36706 64932 38220
rect 64988 38162 65044 38220
rect 64988 38110 64990 38162
rect 65042 38110 65044 38162
rect 64988 38098 65044 38110
rect 64876 36654 64878 36706
rect 64930 36654 64932 36706
rect 64876 36642 64932 36654
rect 64988 37380 65044 37390
rect 64988 36594 65044 37324
rect 65212 37380 65268 40348
rect 65324 40338 65380 40348
rect 65548 41076 65604 41086
rect 65548 38834 65604 41020
rect 65548 38782 65550 38834
rect 65602 38782 65604 38834
rect 65548 38612 65604 38782
rect 65324 38556 65604 38612
rect 65660 38724 65716 41244
rect 65996 41188 66052 41198
rect 65996 41094 66052 41132
rect 66444 41188 66500 42478
rect 67116 41860 67172 41870
rect 67116 41858 67396 41860
rect 67116 41806 67118 41858
rect 67170 41806 67396 41858
rect 67116 41804 67396 41806
rect 67116 41794 67172 41804
rect 66444 41122 66500 41132
rect 67340 41074 67396 41804
rect 67340 41022 67342 41074
rect 67394 41022 67396 41074
rect 67340 41010 67396 41022
rect 67452 40402 67508 45052
rect 67452 40350 67454 40402
rect 67506 40350 67508 40402
rect 67452 40338 67508 40350
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65324 38052 65380 38556
rect 65548 38164 65604 38174
rect 65660 38164 65716 38668
rect 66220 38722 66276 38734
rect 66220 38670 66222 38722
rect 66274 38670 66276 38722
rect 66220 38668 66276 38670
rect 67564 38668 67620 46284
rect 68124 45890 68180 46508
rect 68124 45838 68126 45890
rect 68178 45838 68180 45890
rect 68124 45826 68180 45838
rect 68236 45668 68292 47182
rect 68348 45778 68404 47292
rect 68460 47346 68516 48188
rect 68684 47908 68740 48188
rect 68684 47842 68740 47852
rect 69244 47684 69300 50372
rect 69468 50370 69748 50372
rect 69468 50318 69694 50370
rect 69746 50318 69748 50370
rect 69468 50316 69748 50318
rect 69356 49922 69412 49934
rect 69356 49870 69358 49922
rect 69410 49870 69412 49922
rect 69356 48020 69412 49870
rect 69468 48354 69524 50316
rect 69692 50306 69748 50316
rect 69692 49812 69748 49822
rect 69692 49718 69748 49756
rect 69580 49028 69636 49038
rect 69580 48934 69636 48972
rect 69468 48302 69470 48354
rect 69522 48302 69524 48354
rect 69468 48290 69524 48302
rect 69356 47954 69412 47964
rect 69244 47628 69524 47684
rect 68460 47294 68462 47346
rect 68514 47294 68516 47346
rect 68460 47282 68516 47294
rect 68572 47348 68628 47358
rect 68572 47254 68628 47292
rect 69468 47346 69524 47628
rect 69580 47460 69636 47470
rect 69580 47366 69636 47404
rect 69468 47294 69470 47346
rect 69522 47294 69524 47346
rect 69244 47234 69300 47246
rect 69244 47182 69246 47234
rect 69298 47182 69300 47234
rect 68460 47124 68516 47134
rect 68460 45890 68516 47068
rect 69244 47124 69300 47182
rect 69244 47058 69300 47068
rect 69468 46564 69524 47294
rect 69692 46564 69748 46574
rect 69468 46508 69692 46564
rect 69692 46432 69748 46508
rect 69804 46116 69860 50540
rect 70364 50540 70532 50596
rect 70700 51266 70756 51278
rect 70700 51214 70702 51266
rect 70754 51214 70756 51266
rect 70700 50596 70756 51214
rect 71036 51268 71092 51278
rect 71708 51268 71764 51278
rect 71036 51266 71764 51268
rect 71036 51214 71038 51266
rect 71090 51214 71710 51266
rect 71762 51214 71764 51266
rect 71036 51212 71764 51214
rect 71036 51202 71092 51212
rect 70028 50482 70084 50494
rect 70028 50430 70030 50482
rect 70082 50430 70084 50482
rect 69916 50370 69972 50382
rect 69916 50318 69918 50370
rect 69970 50318 69972 50370
rect 69916 49252 69972 50318
rect 70028 50036 70084 50430
rect 70364 50428 70420 50540
rect 70700 50530 70756 50540
rect 71148 50596 71204 50606
rect 71148 50502 71204 50540
rect 70028 49970 70084 49980
rect 70252 50372 70420 50428
rect 70476 50372 70532 50382
rect 69916 49186 69972 49196
rect 70252 47572 70308 50372
rect 70364 49812 70420 49822
rect 70476 49812 70532 50316
rect 70420 49756 70532 49812
rect 70588 49922 70644 49934
rect 70588 49870 70590 49922
rect 70642 49870 70644 49922
rect 70364 49680 70420 49756
rect 70588 49476 70644 49870
rect 71260 49810 71316 51212
rect 71708 50372 71764 51212
rect 71708 50306 71764 50316
rect 71820 50482 71876 50494
rect 71820 50430 71822 50482
rect 71874 50430 71876 50482
rect 71820 50036 71876 50430
rect 71932 50036 71988 50046
rect 71820 50034 71988 50036
rect 71820 49982 71934 50034
rect 71986 49982 71988 50034
rect 71820 49980 71988 49982
rect 71932 49970 71988 49980
rect 72156 50036 72212 50046
rect 71260 49758 71262 49810
rect 71314 49758 71316 49810
rect 71260 49746 71316 49758
rect 71484 49922 71540 49934
rect 71484 49870 71486 49922
rect 71538 49870 71540 49922
rect 70588 49410 70644 49420
rect 70812 49476 70868 49486
rect 70252 47516 70532 47572
rect 70028 47348 70084 47358
rect 70028 47254 70084 47292
rect 70364 47346 70420 47358
rect 70364 47294 70366 47346
rect 70418 47294 70420 47346
rect 70252 47234 70308 47246
rect 70252 47182 70254 47234
rect 70306 47182 70308 47234
rect 70140 46564 70196 46574
rect 70140 46470 70196 46508
rect 68460 45838 68462 45890
rect 68514 45838 68516 45890
rect 68460 45826 68516 45838
rect 69692 46060 69860 46116
rect 68348 45726 68350 45778
rect 68402 45726 68404 45778
rect 68348 45714 68404 45726
rect 67676 45612 68292 45668
rect 67676 45218 67732 45612
rect 67676 45166 67678 45218
rect 67730 45166 67732 45218
rect 67676 45154 67732 45166
rect 69468 45108 69524 45118
rect 69468 44322 69524 45052
rect 69468 44270 69470 44322
rect 69522 44270 69524 44322
rect 69468 44258 69524 44270
rect 68012 43876 68068 43886
rect 67676 41188 67732 41198
rect 67676 41094 67732 41132
rect 66220 38612 66500 38668
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 66444 38276 66500 38612
rect 65548 38162 65716 38164
rect 65548 38110 65550 38162
rect 65602 38110 65716 38162
rect 65548 38108 65716 38110
rect 66220 38220 66500 38276
rect 67452 38612 67620 38668
rect 65548 38098 65604 38108
rect 65324 37492 65380 37996
rect 66220 37938 66276 38220
rect 66220 37886 66222 37938
rect 66274 37886 66276 37938
rect 66220 37874 66276 37886
rect 66556 37940 66612 37950
rect 66556 37846 66612 37884
rect 67228 37940 67284 37950
rect 67452 37940 67508 38612
rect 67564 38052 67620 38062
rect 67564 37958 67620 37996
rect 67228 37846 67284 37884
rect 67340 37884 67508 37940
rect 65772 37492 65828 37502
rect 65324 37490 65828 37492
rect 65324 37438 65326 37490
rect 65378 37438 65774 37490
rect 65826 37438 65828 37490
rect 65324 37436 65828 37438
rect 65324 37426 65380 37436
rect 65772 37426 65828 37436
rect 65212 37314 65268 37324
rect 66780 37268 66836 37278
rect 66332 37212 66780 37268
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 64988 36542 64990 36594
rect 65042 36542 65044 36594
rect 64988 36530 65044 36542
rect 65436 36706 65492 36718
rect 65436 36654 65438 36706
rect 65490 36654 65492 36706
rect 65436 36594 65492 36654
rect 65436 36542 65438 36594
rect 65490 36542 65492 36594
rect 65436 36530 65492 36542
rect 64540 35870 64542 35922
rect 64594 35870 64596 35922
rect 64540 35858 64596 35870
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 64316 34974 64318 35026
rect 64370 34974 64372 35026
rect 64316 34962 64372 34974
rect 66108 35028 66164 35038
rect 63868 34916 63924 34926
rect 63868 34020 63924 34860
rect 65324 34916 65380 34926
rect 65324 34822 65380 34860
rect 66108 34914 66164 34972
rect 66108 34862 66110 34914
rect 66162 34862 66164 34914
rect 66108 34850 66164 34862
rect 65884 34802 65940 34814
rect 65884 34750 65886 34802
rect 65938 34750 65940 34802
rect 64988 34690 65044 34702
rect 64988 34638 64990 34690
rect 65042 34638 65044 34690
rect 64540 34356 64596 34366
rect 64540 34262 64596 34300
rect 64988 34244 65044 34638
rect 65884 34356 65940 34750
rect 65884 34290 65940 34300
rect 66220 34356 66276 34366
rect 66332 34356 66388 37212
rect 66780 37174 66836 37212
rect 67340 36932 67396 37884
rect 68012 37268 68068 43820
rect 69356 43428 69412 43438
rect 69356 43334 69412 43372
rect 68572 42868 68628 42878
rect 68572 42774 68628 42812
rect 69356 42868 69412 42878
rect 69356 42754 69412 42812
rect 69356 42702 69358 42754
rect 69410 42702 69412 42754
rect 69356 42690 69412 42702
rect 68684 41860 68740 41870
rect 68684 41298 68740 41804
rect 69244 41860 69300 41870
rect 69244 41766 69300 41804
rect 69692 41636 69748 46060
rect 70252 46004 70308 47182
rect 70364 47236 70420 47294
rect 70364 47170 70420 47180
rect 69804 45948 70308 46004
rect 69804 44994 69860 45948
rect 70140 45666 70196 45678
rect 70140 45614 70142 45666
rect 70194 45614 70196 45666
rect 70140 45108 70196 45614
rect 70140 45042 70196 45052
rect 69804 44942 69806 44994
rect 69858 44942 69860 44994
rect 69804 44930 69860 44942
rect 70364 44994 70420 45006
rect 70364 44942 70366 44994
rect 70418 44942 70420 44994
rect 70252 44210 70308 44222
rect 70252 44158 70254 44210
rect 70306 44158 70308 44210
rect 70252 43762 70308 44158
rect 70252 43710 70254 43762
rect 70306 43710 70308 43762
rect 70252 43698 70308 43710
rect 70028 43540 70084 43550
rect 70028 43446 70084 43484
rect 70364 43428 70420 44942
rect 70364 43362 70420 43372
rect 70476 42084 70532 47516
rect 70812 47570 70868 49420
rect 71484 49364 71540 49870
rect 71484 49298 71540 49308
rect 71932 49364 71988 49374
rect 70812 47518 70814 47570
rect 70866 47518 70868 47570
rect 70812 47460 70868 47518
rect 70812 47394 70868 47404
rect 71260 48692 71316 48702
rect 71260 47236 71316 48636
rect 71596 48356 71652 48366
rect 71596 48130 71652 48300
rect 71596 48078 71598 48130
rect 71650 48078 71652 48130
rect 71596 48066 71652 48078
rect 71260 47142 71316 47180
rect 71932 47460 71988 49308
rect 72044 48468 72100 48478
rect 72156 48468 72212 49980
rect 72268 49922 72324 51324
rect 72268 49870 72270 49922
rect 72322 49870 72324 49922
rect 72268 49858 72324 49870
rect 72492 50148 72548 50158
rect 72044 48466 72212 48468
rect 72044 48414 72046 48466
rect 72098 48414 72212 48466
rect 72044 48412 72212 48414
rect 72380 48468 72436 48478
rect 72044 48402 72100 48412
rect 72268 48356 72324 48366
rect 72268 48262 72324 48300
rect 72380 48354 72436 48412
rect 72380 48302 72382 48354
rect 72434 48302 72436 48354
rect 72380 48290 72436 48302
rect 72156 47460 72212 47470
rect 72492 47460 72548 50092
rect 71932 47458 72212 47460
rect 71932 47406 72158 47458
rect 72210 47406 72212 47458
rect 71932 47404 72212 47406
rect 70588 46900 70644 46910
rect 70588 46806 70644 46844
rect 71932 46898 71988 47404
rect 72156 47394 72212 47404
rect 72380 47404 72548 47460
rect 72268 47348 72324 47358
rect 72268 47254 72324 47292
rect 71932 46846 71934 46898
rect 71986 46846 71988 46898
rect 71932 46834 71988 46846
rect 70924 45332 70980 45342
rect 71372 45332 71428 45342
rect 72380 45332 72436 47404
rect 72492 47234 72548 47246
rect 72492 47182 72494 47234
rect 72546 47182 72548 47234
rect 72492 46788 72548 47182
rect 72492 46722 72548 46732
rect 70924 45330 72436 45332
rect 70924 45278 70926 45330
rect 70978 45278 71374 45330
rect 71426 45278 72436 45330
rect 70924 45276 72436 45278
rect 70924 45266 70980 45276
rect 71372 45266 71428 45276
rect 71260 44436 71316 44446
rect 70924 43540 70980 43550
rect 70924 43446 70980 43484
rect 71260 43538 71316 44380
rect 71260 43486 71262 43538
rect 71314 43486 71316 43538
rect 71260 43474 71316 43486
rect 71484 43650 71540 43662
rect 71484 43598 71486 43650
rect 71538 43598 71540 43650
rect 71484 43428 71540 43598
rect 71484 43362 71540 43372
rect 71708 42194 71764 45276
rect 72268 45108 72324 45118
rect 72268 44100 72324 45052
rect 72044 43652 72100 43662
rect 72044 43558 72100 43596
rect 71708 42142 71710 42194
rect 71762 42142 71764 42194
rect 70812 42084 70868 42094
rect 70476 42082 70868 42084
rect 70476 42030 70814 42082
rect 70866 42030 70868 42082
rect 70476 42028 70868 42030
rect 70476 41860 70532 42028
rect 70812 42018 70868 42028
rect 70924 41970 70980 41982
rect 70924 41918 70926 41970
rect 70978 41918 70980 41970
rect 70476 41794 70532 41804
rect 70812 41860 70868 41870
rect 69916 41746 69972 41758
rect 69916 41694 69918 41746
rect 69970 41694 69972 41746
rect 69692 41580 69860 41636
rect 68684 41246 68686 41298
rect 68738 41246 68740 41298
rect 68684 41234 68740 41246
rect 69468 41300 69524 41310
rect 69468 41206 69524 41244
rect 68124 40290 68180 40302
rect 68124 40238 68126 40290
rect 68178 40238 68180 40290
rect 68124 39508 68180 40238
rect 69692 39620 69748 39630
rect 69244 39618 69748 39620
rect 69244 39566 69694 39618
rect 69746 39566 69748 39618
rect 69244 39564 69748 39566
rect 68236 39508 68292 39518
rect 68124 39506 68292 39508
rect 68124 39454 68238 39506
rect 68290 39454 68292 39506
rect 68124 39452 68292 39454
rect 68236 39442 68292 39452
rect 68572 39506 68628 39518
rect 68572 39454 68574 39506
rect 68626 39454 68628 39506
rect 68572 39060 68628 39454
rect 68572 38994 68628 39004
rect 68236 38724 68292 38734
rect 68348 38724 68404 38734
rect 68292 38722 68404 38724
rect 68292 38670 68350 38722
rect 68402 38670 68404 38722
rect 68292 38668 68404 38670
rect 68236 37938 68292 38668
rect 68348 38658 68404 38668
rect 68236 37886 68238 37938
rect 68290 37886 68292 37938
rect 68236 37874 68292 37886
rect 68348 38164 68404 38174
rect 68348 38050 68404 38108
rect 68348 37998 68350 38050
rect 68402 37998 68404 38050
rect 69244 38164 69300 39564
rect 69692 39554 69748 39564
rect 69692 39060 69748 39070
rect 69692 38966 69748 39004
rect 69804 38724 69860 41580
rect 69916 41188 69972 41694
rect 69916 41122 69972 41132
rect 70252 41746 70308 41758
rect 70252 41694 70254 41746
rect 70306 41694 70308 41746
rect 69916 40964 69972 40974
rect 69916 40870 69972 40908
rect 70252 40292 70308 41694
rect 70700 41636 70756 41646
rect 70364 41300 70420 41310
rect 70364 41206 70420 41244
rect 70700 40626 70756 41580
rect 70812 41298 70868 41804
rect 70812 41246 70814 41298
rect 70866 41246 70868 41298
rect 70812 40964 70868 41246
rect 70924 41300 70980 41918
rect 71708 41972 71764 42142
rect 71708 41906 71764 41916
rect 72268 42866 72324 44044
rect 72380 44436 72436 44446
rect 72380 43764 72436 44380
rect 72380 43698 72436 43708
rect 72268 42814 72270 42866
rect 72322 42814 72324 42866
rect 72156 41860 72212 41870
rect 72044 41858 72212 41860
rect 72044 41806 72158 41858
rect 72210 41806 72212 41858
rect 72044 41804 72212 41806
rect 72044 41748 72100 41804
rect 72156 41794 72212 41804
rect 70924 41234 70980 41244
rect 71932 41692 72100 41748
rect 70812 40898 70868 40908
rect 71260 41188 71316 41198
rect 70700 40574 70702 40626
rect 70754 40574 70756 40626
rect 70700 40562 70756 40574
rect 71260 40626 71316 41132
rect 71820 41188 71876 41198
rect 71820 41094 71876 41132
rect 71260 40574 71262 40626
rect 71314 40574 71316 40626
rect 70028 40290 70308 40292
rect 70028 40238 70254 40290
rect 70306 40238 70308 40290
rect 70028 40236 70308 40238
rect 70028 38834 70084 40236
rect 70252 40226 70308 40236
rect 70252 39732 70308 39742
rect 70252 39618 70308 39676
rect 70700 39732 70756 39742
rect 70700 39638 70756 39676
rect 71260 39732 71316 40574
rect 71260 39666 71316 39676
rect 71708 40290 71764 40302
rect 71708 40238 71710 40290
rect 71762 40238 71764 40290
rect 70252 39566 70254 39618
rect 70306 39566 70308 39618
rect 70252 39554 70308 39566
rect 70028 38782 70030 38834
rect 70082 38782 70084 38834
rect 70028 38770 70084 38782
rect 70700 39060 70756 39070
rect 70700 38834 70756 39004
rect 71372 39060 71428 39070
rect 71372 38966 71428 39004
rect 70700 38782 70702 38834
rect 70754 38782 70756 38834
rect 70700 38770 70756 38782
rect 70812 38946 70868 38958
rect 70812 38894 70814 38946
rect 70866 38894 70868 38946
rect 69244 38032 69300 38108
rect 69692 38164 69748 38174
rect 69804 38164 69860 38668
rect 69692 38162 69860 38164
rect 69692 38110 69694 38162
rect 69746 38110 69860 38162
rect 69692 38108 69860 38110
rect 69692 38098 69748 38108
rect 69580 38052 69636 38062
rect 68348 37716 68404 37998
rect 68348 37650 68404 37660
rect 68012 37212 68292 37268
rect 67452 37156 67508 37166
rect 67452 37154 68068 37156
rect 67452 37102 67454 37154
rect 67506 37102 68068 37154
rect 67452 37100 68068 37102
rect 67452 37090 67508 37100
rect 67340 36876 67508 36932
rect 66668 35588 66724 35598
rect 66668 35494 66724 35532
rect 67228 35588 67284 35598
rect 66668 35028 66724 35038
rect 66668 34934 66724 34972
rect 66220 34354 66388 34356
rect 66220 34302 66222 34354
rect 66274 34302 66388 34354
rect 66220 34300 66388 34302
rect 66220 34290 66276 34300
rect 65436 34244 65492 34254
rect 64988 34178 65044 34188
rect 65100 34242 65492 34244
rect 65100 34190 65438 34242
rect 65490 34190 65492 34242
rect 65100 34188 65492 34190
rect 63868 33926 63924 33964
rect 65100 33796 65156 34188
rect 65436 34178 65492 34188
rect 65772 34244 65828 34254
rect 65772 34150 65828 34188
rect 64204 33740 65156 33796
rect 65916 33740 66180 33750
rect 64204 33458 64260 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 64204 33406 64206 33458
rect 64258 33406 64260 33458
rect 64204 33394 64260 33406
rect 64988 33348 65044 33358
rect 64988 33254 65044 33292
rect 65772 33348 65828 33358
rect 62860 32786 63700 32788
rect 62860 32734 63534 32786
rect 63586 32734 63700 32786
rect 62860 32732 63700 32734
rect 62636 32676 62692 32686
rect 62636 32582 62692 32620
rect 62076 32564 62132 32574
rect 61964 32562 62132 32564
rect 61964 32510 62078 32562
rect 62130 32510 62132 32562
rect 61964 32508 62132 32510
rect 62076 32498 62132 32508
rect 62860 32562 62916 32732
rect 63532 32722 63588 32732
rect 62860 32510 62862 32562
rect 62914 32510 62916 32562
rect 62860 32498 62916 32510
rect 65772 32562 65828 33292
rect 66332 33348 66388 34300
rect 67228 34130 67284 35532
rect 67228 34078 67230 34130
rect 67282 34078 67284 34130
rect 67228 34066 67284 34078
rect 67340 34690 67396 34702
rect 67340 34638 67342 34690
rect 67394 34638 67396 34690
rect 66332 33282 66388 33292
rect 66444 33236 66500 33246
rect 67340 33236 67396 34638
rect 66444 33234 66724 33236
rect 66444 33182 66446 33234
rect 66498 33182 66724 33234
rect 66444 33180 66724 33182
rect 66444 33170 66500 33180
rect 65772 32510 65774 32562
rect 65826 32510 65828 32562
rect 65772 32498 65828 32510
rect 66444 32450 66500 32462
rect 66444 32398 66446 32450
rect 66498 32398 66500 32450
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 61404 31838 61406 31890
rect 61458 31838 61460 31890
rect 61404 31826 61460 31838
rect 66444 31668 66500 32398
rect 66444 31602 66500 31612
rect 66668 31666 66724 33180
rect 67004 33180 67396 33236
rect 67004 31778 67060 33180
rect 67004 31726 67006 31778
rect 67058 31726 67060 31778
rect 67004 31714 67060 31726
rect 67452 31780 67508 36876
rect 68012 36370 68068 37100
rect 68012 36318 68014 36370
rect 68066 36318 68068 36370
rect 68012 36306 68068 36318
rect 67676 34914 67732 34926
rect 67676 34862 67678 34914
rect 67730 34862 67732 34914
rect 67676 32452 67732 34862
rect 68236 34916 68292 37212
rect 69580 37156 69636 37996
rect 70140 37268 70196 37278
rect 69580 37154 69860 37156
rect 69580 37102 69582 37154
rect 69634 37102 69860 37154
rect 69580 37100 69860 37102
rect 69580 37090 69636 37100
rect 69804 36706 69860 37100
rect 69804 36654 69806 36706
rect 69858 36654 69860 36706
rect 69804 36642 69860 36654
rect 70140 37154 70196 37212
rect 70140 37102 70142 37154
rect 70194 37102 70196 37154
rect 68348 36372 68404 36382
rect 68348 36278 68404 36316
rect 69468 36372 69524 36382
rect 69468 36278 69524 36316
rect 68236 34802 68292 34860
rect 68236 34750 68238 34802
rect 68290 34750 68292 34802
rect 68236 34738 68292 34750
rect 68460 34914 68516 34926
rect 68460 34862 68462 34914
rect 68514 34862 68516 34914
rect 68460 34692 68516 34862
rect 68460 34626 68516 34636
rect 68572 34916 68628 34926
rect 68572 33458 68628 34860
rect 69692 34916 69748 34926
rect 69692 34822 69748 34860
rect 69356 34692 69412 34702
rect 69356 34598 69412 34636
rect 70140 34242 70196 37102
rect 70588 36820 70644 36830
rect 70588 36482 70644 36764
rect 70588 36430 70590 36482
rect 70642 36430 70644 36482
rect 70588 36418 70644 36430
rect 70364 36372 70420 36382
rect 70140 34190 70142 34242
rect 70194 34190 70196 34242
rect 70140 34178 70196 34190
rect 70252 36316 70364 36372
rect 68572 33406 68574 33458
rect 68626 33406 68628 33458
rect 68572 33394 68628 33406
rect 68684 33348 68740 33358
rect 67676 32386 67732 32396
rect 68572 32452 68628 32462
rect 68572 32358 68628 32396
rect 67452 31714 67508 31724
rect 68012 32340 68068 32350
rect 68012 31778 68068 32284
rect 68572 31892 68628 31902
rect 68684 31892 68740 33292
rect 69692 33348 69748 33358
rect 69692 33254 69748 33292
rect 70252 33124 70308 36316
rect 70364 36240 70420 36316
rect 70812 36372 70868 38894
rect 71148 36820 71204 36830
rect 71148 36594 71204 36764
rect 71708 36820 71764 40238
rect 71932 39060 71988 41692
rect 72268 41636 72324 42814
rect 72044 41580 72268 41636
rect 72044 40404 72100 41580
rect 72268 41570 72324 41580
rect 72268 41412 72324 41422
rect 72268 41298 72324 41356
rect 72268 41246 72270 41298
rect 72322 41246 72324 41298
rect 72268 41234 72324 41246
rect 72268 41076 72324 41086
rect 72268 40626 72324 41020
rect 72268 40574 72270 40626
rect 72322 40574 72324 40626
rect 72268 40562 72324 40574
rect 72044 39618 72100 40348
rect 72044 39566 72046 39618
rect 72098 39566 72100 39618
rect 72044 39554 72100 39566
rect 71932 38994 71988 39004
rect 71708 36754 71764 36764
rect 71820 38722 71876 38734
rect 71820 38670 71822 38722
rect 71874 38670 71876 38722
rect 71148 36542 71150 36594
rect 71202 36542 71204 36594
rect 71148 36530 71204 36542
rect 70812 36306 70868 36316
rect 71596 36372 71652 36382
rect 71820 36372 71876 38670
rect 72604 38668 72660 52108
rect 72828 52098 72884 52108
rect 72716 48468 72772 48478
rect 72716 46898 72772 48412
rect 72716 46846 72718 46898
rect 72770 46846 72772 46898
rect 72716 46834 72772 46846
rect 72828 47348 72884 47358
rect 72940 47348 72996 53340
rect 73052 52836 73108 53454
rect 73276 53172 73332 58270
rect 73388 57876 73444 59836
rect 73500 59332 73556 60732
rect 73724 59556 73780 61516
rect 73948 61506 74004 61516
rect 73948 60002 74004 60014
rect 73948 59950 73950 60002
rect 74002 59950 74004 60002
rect 73948 59780 74004 59950
rect 74060 59892 74116 62188
rect 74172 64204 74340 64260
rect 74172 61794 74228 64204
rect 74396 64146 74452 64158
rect 74396 64094 74398 64146
rect 74450 64094 74452 64146
rect 74396 62804 74452 64094
rect 74732 63028 74788 66108
rect 74956 66164 75012 66174
rect 74956 66070 75012 66108
rect 74956 65490 75012 65502
rect 74956 65438 74958 65490
rect 75010 65438 75012 65490
rect 74956 64708 75012 65438
rect 74956 64642 75012 64652
rect 74956 63924 75012 63934
rect 74732 62972 74900 63028
rect 74396 62738 74452 62748
rect 74732 62804 74788 62814
rect 74508 62468 74564 62478
rect 74396 62020 74452 62030
rect 74172 61742 74174 61794
rect 74226 61742 74228 61794
rect 74172 61730 74228 61742
rect 74284 61908 74340 61918
rect 74284 61682 74340 61852
rect 74284 61630 74286 61682
rect 74338 61630 74340 61682
rect 74284 61618 74340 61630
rect 74396 61570 74452 61964
rect 74396 61518 74398 61570
rect 74450 61518 74452 61570
rect 74396 61506 74452 61518
rect 74508 60228 74564 62412
rect 74508 60172 74676 60228
rect 74508 60004 74564 60014
rect 74508 59910 74564 59948
rect 74060 59890 74228 59892
rect 74060 59838 74062 59890
rect 74114 59838 74228 59890
rect 74060 59836 74228 59838
rect 74060 59826 74116 59836
rect 73724 59490 73780 59500
rect 73892 59724 74004 59780
rect 73500 59266 73556 59276
rect 73892 58996 73948 59724
rect 73836 58940 73948 58996
rect 73836 58660 73892 58940
rect 73500 58604 73892 58660
rect 73500 58434 73556 58604
rect 73500 58382 73502 58434
rect 73554 58382 73556 58434
rect 73500 58100 73556 58382
rect 73612 58436 73668 58446
rect 73612 58322 73668 58380
rect 73612 58270 73614 58322
rect 73666 58270 73668 58322
rect 73612 58258 73668 58270
rect 74060 58434 74116 58446
rect 74060 58382 74062 58434
rect 74114 58382 74116 58434
rect 74060 58324 74116 58382
rect 74172 58436 74228 59836
rect 74396 59330 74452 59342
rect 74396 59278 74398 59330
rect 74450 59278 74452 59330
rect 74172 58370 74228 58380
rect 74284 58548 74340 58558
rect 74060 58100 74116 58268
rect 73500 58044 73668 58100
rect 73500 57876 73556 57886
rect 73388 57874 73556 57876
rect 73388 57822 73502 57874
rect 73554 57822 73556 57874
rect 73388 57820 73556 57822
rect 73388 57652 73444 57820
rect 73500 57810 73556 57820
rect 73388 57586 73444 57596
rect 73612 57762 73668 58044
rect 74060 58034 74116 58044
rect 73612 57710 73614 57762
rect 73666 57710 73668 57762
rect 73500 57428 73556 57438
rect 73388 57426 73556 57428
rect 73388 57374 73502 57426
rect 73554 57374 73556 57426
rect 73388 57372 73556 57374
rect 73388 55412 73444 57372
rect 73500 57362 73556 57372
rect 73612 56978 73668 57710
rect 74172 57876 74228 57886
rect 73612 56926 73614 56978
rect 73666 56926 73668 56978
rect 73612 56914 73668 56926
rect 73724 57652 73780 57662
rect 73724 56306 73780 57596
rect 74060 57426 74116 57438
rect 74060 57374 74062 57426
rect 74114 57374 74116 57426
rect 74060 56980 74116 57374
rect 74060 56914 74116 56924
rect 73724 56254 73726 56306
rect 73778 56254 73780 56306
rect 73724 56242 73780 56254
rect 73836 56866 73892 56878
rect 73836 56814 73838 56866
rect 73890 56814 73892 56866
rect 73500 56196 73556 56206
rect 73500 56102 73556 56140
rect 73836 56196 73892 56814
rect 74172 56866 74228 57820
rect 74284 57652 74340 58492
rect 74396 58436 74452 59278
rect 74620 58996 74676 60172
rect 74620 58930 74676 58940
rect 74620 58436 74676 58446
rect 74396 58434 74676 58436
rect 74396 58382 74622 58434
rect 74674 58382 74676 58434
rect 74396 58380 74676 58382
rect 74620 58324 74676 58380
rect 74620 58258 74676 58268
rect 74732 57876 74788 62748
rect 74844 62468 74900 62972
rect 74844 62402 74900 62412
rect 74956 61572 75012 63868
rect 75068 63922 75124 67564
rect 75068 63870 75070 63922
rect 75122 63870 75124 63922
rect 75068 63858 75124 63870
rect 75180 63700 75236 68348
rect 75292 67732 75348 68572
rect 75292 67666 75348 67676
rect 75516 67956 75572 67966
rect 75404 67620 75460 67630
rect 75404 67526 75460 67564
rect 75516 67284 75572 67900
rect 75516 67218 75572 67228
rect 75740 67956 75796 67966
rect 76188 67956 76244 69132
rect 76300 69122 76356 69132
rect 76300 68628 76356 68638
rect 76300 68534 76356 68572
rect 75740 67954 76244 67956
rect 75740 67902 75742 67954
rect 75794 67902 76190 67954
rect 76242 67902 76244 67954
rect 75740 67900 76244 67902
rect 75740 67172 75796 67900
rect 76188 67890 76244 67900
rect 76412 67508 76468 70702
rect 75740 67106 75796 67116
rect 75964 67452 76468 67508
rect 75964 67170 76020 67452
rect 76076 67284 76132 67294
rect 76076 67282 76244 67284
rect 76076 67230 76078 67282
rect 76130 67230 76244 67282
rect 76076 67228 76244 67230
rect 76076 67218 76132 67228
rect 75964 67118 75966 67170
rect 76018 67118 76020 67170
rect 75404 66946 75460 66958
rect 75404 66894 75406 66946
rect 75458 66894 75460 66946
rect 75404 65380 75460 66894
rect 75516 66948 75572 66958
rect 75516 66274 75572 66892
rect 75516 66222 75518 66274
rect 75570 66222 75572 66274
rect 75516 66210 75572 66222
rect 75964 66388 76020 67118
rect 75852 66164 75908 66174
rect 75964 66164 76020 66332
rect 75852 66162 76020 66164
rect 75852 66110 75854 66162
rect 75906 66110 76020 66162
rect 75852 66108 76020 66110
rect 76076 66834 76132 66846
rect 76076 66782 76078 66834
rect 76130 66782 76132 66834
rect 75852 66098 75908 66108
rect 75404 63924 75460 65324
rect 75404 63858 75460 63868
rect 75740 65940 75796 65950
rect 75180 63634 75236 63644
rect 75740 63700 75796 65884
rect 75964 65602 76020 65614
rect 75964 65550 75966 65602
rect 76018 65550 76020 65602
rect 75740 63634 75796 63644
rect 75852 64594 75908 64606
rect 75852 64542 75854 64594
rect 75906 64542 75908 64594
rect 75404 63588 75460 63598
rect 75404 62578 75460 63532
rect 75404 62526 75406 62578
rect 75458 62526 75460 62578
rect 75404 62514 75460 62526
rect 75516 63476 75572 63486
rect 75404 62356 75460 62394
rect 75404 62290 75460 62300
rect 75404 62132 75460 62142
rect 75404 61684 75460 62076
rect 75180 61572 75236 61582
rect 74956 61570 75236 61572
rect 74956 61518 75182 61570
rect 75234 61518 75236 61570
rect 74956 61516 75236 61518
rect 75180 61506 75236 61516
rect 75404 61570 75460 61628
rect 75404 61518 75406 61570
rect 75458 61518 75460 61570
rect 75404 61506 75460 61518
rect 75180 61348 75236 61358
rect 74956 60226 75012 60238
rect 74956 60174 74958 60226
rect 75010 60174 75012 60226
rect 74284 57520 74340 57596
rect 74396 57820 74788 57876
rect 74844 59444 74900 59454
rect 74172 56814 74174 56866
rect 74226 56814 74228 56866
rect 74172 56644 74228 56814
rect 74172 56578 74228 56588
rect 73948 56308 74004 56318
rect 74396 56308 74452 57820
rect 74844 57762 74900 59388
rect 74844 57710 74846 57762
rect 74898 57710 74900 57762
rect 74844 57698 74900 57710
rect 74732 57650 74788 57662
rect 74732 57598 74734 57650
rect 74786 57598 74788 57650
rect 74732 57092 74788 57598
rect 74956 57204 75012 60174
rect 75068 57764 75124 57774
rect 75068 57650 75124 57708
rect 75068 57598 75070 57650
rect 75122 57598 75124 57650
rect 75068 57586 75124 57598
rect 74956 57138 75012 57148
rect 74732 57026 74788 57036
rect 73948 56214 74004 56252
rect 74284 56252 74452 56308
rect 74844 56980 74900 56990
rect 73388 55346 73444 55356
rect 73388 55186 73444 55198
rect 73388 55134 73390 55186
rect 73442 55134 73444 55186
rect 73388 54404 73444 55134
rect 73836 54514 73892 56140
rect 74060 55860 74116 55870
rect 74060 55858 74228 55860
rect 74060 55806 74062 55858
rect 74114 55806 74228 55858
rect 74060 55804 74228 55806
rect 74060 55794 74116 55804
rect 73836 54462 73838 54514
rect 73890 54462 73892 54514
rect 73836 54450 73892 54462
rect 74060 54740 74116 54750
rect 74060 54514 74116 54684
rect 74060 54462 74062 54514
rect 74114 54462 74116 54514
rect 74060 54450 74116 54462
rect 73388 54402 73556 54404
rect 73388 54350 73390 54402
rect 73442 54350 73556 54402
rect 73388 54348 73556 54350
rect 73388 54338 73444 54348
rect 73500 53620 73556 54348
rect 73612 54290 73668 54302
rect 73612 54238 73614 54290
rect 73666 54238 73668 54290
rect 73612 53954 73668 54238
rect 73612 53902 73614 53954
rect 73666 53902 73668 53954
rect 73612 53890 73668 53902
rect 73500 53508 73556 53564
rect 73500 53506 73780 53508
rect 73500 53454 73502 53506
rect 73554 53454 73780 53506
rect 73500 53452 73780 53454
rect 73500 53442 73556 53452
rect 73276 53116 73668 53172
rect 73388 52946 73444 52958
rect 73388 52894 73390 52946
rect 73442 52894 73444 52946
rect 73388 52836 73444 52894
rect 73052 52780 73444 52836
rect 73052 47684 73108 52780
rect 73500 52276 73556 52286
rect 73500 52182 73556 52220
rect 73612 51828 73668 53116
rect 73724 51940 73780 53452
rect 73836 52948 73892 52958
rect 73836 52834 73892 52892
rect 73836 52782 73838 52834
rect 73890 52782 73892 52834
rect 73836 52770 73892 52782
rect 73948 52388 74004 52398
rect 73948 52274 74004 52332
rect 73948 52222 73950 52274
rect 74002 52222 74004 52274
rect 73948 52210 74004 52222
rect 73724 51874 73780 51884
rect 74060 52052 74116 52062
rect 73388 51772 73668 51828
rect 73276 51380 73332 51390
rect 73276 51286 73332 51324
rect 73388 50148 73444 51772
rect 74060 51602 74116 51996
rect 74060 51550 74062 51602
rect 74114 51550 74116 51602
rect 74060 51538 74116 51550
rect 73500 51492 73556 51502
rect 73500 51398 73556 51436
rect 73948 51492 74004 51502
rect 73612 51380 73668 51418
rect 73612 51314 73668 51324
rect 73388 50082 73444 50092
rect 73612 51156 73668 51166
rect 73612 50596 73668 51100
rect 73948 50706 74004 51436
rect 73948 50654 73950 50706
rect 74002 50654 74004 50706
rect 73948 50642 74004 50654
rect 73388 49924 73444 49934
rect 73388 49830 73444 49868
rect 73052 47618 73108 47628
rect 73164 48916 73220 48926
rect 73612 48916 73668 50540
rect 73724 50484 73780 50494
rect 73724 49922 73780 50428
rect 73724 49870 73726 49922
rect 73778 49870 73780 49922
rect 73724 49858 73780 49870
rect 73164 48914 73668 48916
rect 73164 48862 73166 48914
rect 73218 48862 73668 48914
rect 73164 48860 73668 48862
rect 73164 48132 73220 48860
rect 73276 48132 73332 48142
rect 73164 48130 73332 48132
rect 73164 48078 73278 48130
rect 73330 48078 73332 48130
rect 73164 48076 73332 48078
rect 73052 47470 73108 47482
rect 73052 47418 73054 47470
rect 73106 47460 73108 47470
rect 73164 47460 73220 48076
rect 73276 48066 73332 48076
rect 73836 48132 73892 48142
rect 73836 48038 73892 48076
rect 73106 47418 73220 47460
rect 73052 47404 73220 47418
rect 72940 47292 73108 47348
rect 72828 45668 72884 47292
rect 72716 45612 72884 45668
rect 72716 43652 72772 45612
rect 72828 44100 72884 44110
rect 72828 44006 72884 44044
rect 72716 43520 72772 43596
rect 73052 41636 73108 47292
rect 73164 46900 73220 47404
rect 73612 47684 73668 47694
rect 73388 47348 73444 47358
rect 73164 46004 73220 46844
rect 73276 46900 73332 46910
rect 73388 46900 73444 47292
rect 73276 46898 73444 46900
rect 73276 46846 73278 46898
rect 73330 46846 73444 46898
rect 73276 46844 73444 46846
rect 73276 46834 73332 46844
rect 73164 45938 73220 45948
rect 73276 42532 73332 42542
rect 73276 41972 73332 42476
rect 73276 41878 73332 41916
rect 73612 41860 73668 47628
rect 73724 47346 73780 47358
rect 73724 47294 73726 47346
rect 73778 47294 73780 47346
rect 73724 46452 73780 47294
rect 73948 46900 74004 46910
rect 73948 46806 74004 46844
rect 73836 46788 73892 46798
rect 73836 46694 73892 46732
rect 73948 46452 74004 46462
rect 73724 46450 74004 46452
rect 73724 46398 73950 46450
rect 74002 46398 74004 46450
rect 73724 46396 74004 46398
rect 73948 46386 74004 46396
rect 73724 44322 73780 44334
rect 73724 44270 73726 44322
rect 73778 44270 73780 44322
rect 73724 41972 73780 44270
rect 74172 43708 74228 55804
rect 74284 50372 74340 56252
rect 74508 56196 74564 56206
rect 74396 56194 74564 56196
rect 74396 56142 74510 56194
rect 74562 56142 74564 56194
rect 74396 56140 74564 56142
rect 74396 53732 74452 56140
rect 74508 56130 74564 56140
rect 74844 56194 74900 56924
rect 74956 56754 75012 56766
rect 74956 56702 74958 56754
rect 75010 56702 75012 56754
rect 74956 56420 75012 56702
rect 74956 56354 75012 56364
rect 74844 56142 74846 56194
rect 74898 56142 74900 56194
rect 74844 56130 74900 56142
rect 74956 55524 75012 55534
rect 74844 55412 74900 55422
rect 74844 54740 74900 55356
rect 74956 55298 75012 55468
rect 74956 55246 74958 55298
rect 75010 55246 75012 55298
rect 74956 55234 75012 55246
rect 74956 54740 75012 54750
rect 74732 54684 74956 54740
rect 74508 54292 74564 54302
rect 74508 54290 74676 54292
rect 74508 54238 74510 54290
rect 74562 54238 74676 54290
rect 74508 54236 74676 54238
rect 74508 54226 74564 54236
rect 74396 53666 74452 53676
rect 74396 52836 74452 52846
rect 74396 52742 74452 52780
rect 74508 51604 74564 51614
rect 74508 51510 74564 51548
rect 74284 50306 74340 50316
rect 74620 50596 74676 54236
rect 74732 53842 74788 54684
rect 74956 54646 75012 54684
rect 74732 53790 74734 53842
rect 74786 53790 74788 53842
rect 74732 53778 74788 53790
rect 74844 53956 74900 53966
rect 74732 53172 74788 53182
rect 74732 52162 74788 53116
rect 74732 52110 74734 52162
rect 74786 52110 74788 52162
rect 74732 52052 74788 52110
rect 74732 51986 74788 51996
rect 74844 51828 74900 53900
rect 75180 52948 75236 61292
rect 75292 60452 75348 60462
rect 75292 60002 75348 60396
rect 75292 59950 75294 60002
rect 75346 59950 75348 60002
rect 75292 59938 75348 59950
rect 75516 59442 75572 63420
rect 75852 63026 75908 64542
rect 75964 64034 76020 65550
rect 76076 65604 76132 66782
rect 76188 65940 76244 67228
rect 76188 65874 76244 65884
rect 76300 66050 76356 66062
rect 76300 65998 76302 66050
rect 76354 65998 76356 66050
rect 76076 65538 76132 65548
rect 75964 63982 75966 64034
rect 76018 63982 76020 64034
rect 75964 63812 76020 63982
rect 75964 63252 76020 63756
rect 75964 63186 76020 63196
rect 76076 63364 76132 63374
rect 75852 62974 75854 63026
rect 75906 62974 75908 63026
rect 75852 62692 75908 62974
rect 75852 62626 75908 62636
rect 75628 62356 75684 62366
rect 75628 61908 75684 62300
rect 75740 62354 75796 62366
rect 75740 62302 75742 62354
rect 75794 62302 75796 62354
rect 75740 62132 75796 62302
rect 76076 62188 76132 63308
rect 75740 62066 75796 62076
rect 75852 62132 76132 62188
rect 75628 61852 75796 61908
rect 75628 61572 75684 61582
rect 75628 61478 75684 61516
rect 75516 59390 75518 59442
rect 75570 59390 75572 59442
rect 75516 59378 75572 59390
rect 75516 59218 75572 59230
rect 75516 59166 75518 59218
rect 75570 59166 75572 59218
rect 75404 58322 75460 58334
rect 75404 58270 75406 58322
rect 75458 58270 75460 58322
rect 75292 58210 75348 58222
rect 75292 58158 75294 58210
rect 75346 58158 75348 58210
rect 75292 57988 75348 58158
rect 75292 57922 75348 57932
rect 75404 57764 75460 58270
rect 75516 58100 75572 59166
rect 75740 59220 75796 61852
rect 75852 61570 75908 62132
rect 76300 61908 76356 65998
rect 76412 64706 76468 64718
rect 76412 64654 76414 64706
rect 76466 64654 76468 64706
rect 76412 63924 76468 64654
rect 76412 63138 76468 63868
rect 76524 63476 76580 71820
rect 77644 71762 77700 72156
rect 78428 71874 78484 73836
rect 78540 73556 78596 73950
rect 78540 73490 78596 73500
rect 78428 71822 78430 71874
rect 78482 71822 78484 71874
rect 78428 71810 78484 71822
rect 77644 71710 77646 71762
rect 77698 71710 77700 71762
rect 76636 71652 76692 71662
rect 76636 71558 76692 71596
rect 76748 71538 76804 71550
rect 76748 71486 76750 71538
rect 76802 71486 76804 71538
rect 76748 71092 76804 71486
rect 77196 71092 77252 71102
rect 76748 71090 77252 71092
rect 76748 71038 77198 71090
rect 77250 71038 77252 71090
rect 76748 71036 77252 71038
rect 77196 71026 77252 71036
rect 76972 70196 77028 70206
rect 76972 70194 77140 70196
rect 76972 70142 76974 70194
rect 77026 70142 77140 70194
rect 76972 70140 77140 70142
rect 76972 70130 77028 70140
rect 76972 69188 77028 69198
rect 76972 68626 77028 69132
rect 76972 68574 76974 68626
rect 77026 68574 77028 68626
rect 76972 68562 77028 68574
rect 77084 68068 77140 70140
rect 77644 70194 77700 71710
rect 77644 70142 77646 70194
rect 77698 70142 77700 70194
rect 77644 70130 77700 70142
rect 77756 70754 77812 70766
rect 77756 70702 77758 70754
rect 77810 70702 77812 70754
rect 77196 70084 77252 70094
rect 77196 68850 77252 70028
rect 77420 69300 77476 69310
rect 77756 69300 77812 70702
rect 78316 70084 78372 70094
rect 78316 69990 78372 70028
rect 78652 69748 78708 78932
rect 78988 78932 79044 78988
rect 78988 78876 79156 78932
rect 78764 78034 78820 78046
rect 78764 77982 78766 78034
rect 78818 77982 78820 78034
rect 78764 77028 78820 77982
rect 78876 77476 78932 77486
rect 78876 77250 78932 77420
rect 78876 77198 78878 77250
rect 78930 77198 78932 77250
rect 78876 77186 78932 77198
rect 78764 76962 78820 76972
rect 78764 76132 78820 76142
rect 78764 73948 78820 76076
rect 79100 75682 79156 78876
rect 79324 78034 79380 80668
rect 79548 80498 79604 80892
rect 79548 80446 79550 80498
rect 79602 80446 79604 80498
rect 79548 80434 79604 80446
rect 79324 77982 79326 78034
rect 79378 77982 79380 78034
rect 79324 77970 79380 77982
rect 79884 79044 79940 79054
rect 79436 77364 79492 77374
rect 79212 77252 79268 77262
rect 79212 77138 79268 77196
rect 79212 77086 79214 77138
rect 79266 77086 79268 77138
rect 79212 77028 79268 77086
rect 79212 76962 79268 76972
rect 79100 75630 79102 75682
rect 79154 75630 79156 75682
rect 79100 75618 79156 75630
rect 79436 73948 79492 77308
rect 79884 77362 79940 78988
rect 79884 77310 79886 77362
rect 79938 77310 79940 77362
rect 79884 77298 79940 77310
rect 80220 78036 80276 83244
rect 80444 82962 80500 83356
rect 80444 82910 80446 82962
rect 80498 82910 80500 82962
rect 80444 82898 80500 82910
rect 80332 82738 80388 82750
rect 80332 82686 80334 82738
rect 80386 82686 80388 82738
rect 80332 81956 80388 82686
rect 80444 82516 80500 82526
rect 80556 82516 80612 84140
rect 80444 82514 80612 82516
rect 80444 82462 80446 82514
rect 80498 82462 80612 82514
rect 80444 82460 80612 82462
rect 80892 83410 80948 83422
rect 80892 83358 80894 83410
rect 80946 83358 80948 83410
rect 80444 82450 80500 82460
rect 80332 81890 80388 81900
rect 80444 82292 80500 82302
rect 80444 81396 80500 82236
rect 80668 82292 80724 82302
rect 80668 81730 80724 82236
rect 80892 81956 80948 83358
rect 81276 83132 81540 83142
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81276 83066 81540 83076
rect 81452 82626 81508 82638
rect 81452 82574 81454 82626
rect 81506 82574 81508 82626
rect 81452 82292 81508 82574
rect 81452 82226 81508 82236
rect 81116 81956 81172 81966
rect 80892 81954 81172 81956
rect 80892 81902 81118 81954
rect 81170 81902 81172 81954
rect 80892 81900 81172 81902
rect 81116 81890 81172 81900
rect 81452 81956 81508 81966
rect 81676 81956 81732 84364
rect 82012 83412 82068 86828
rect 82348 85764 82404 95788
rect 82908 95778 82964 95788
rect 96636 94892 96900 94902
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96636 94826 96900 94836
rect 96636 93324 96900 93334
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96636 93258 96900 93268
rect 96636 91756 96900 91766
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96636 91690 96900 91700
rect 96636 90188 96900 90198
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96636 90122 96900 90132
rect 90860 89010 90916 89022
rect 90860 88958 90862 89010
rect 90914 88958 90916 89010
rect 87276 87554 87332 87566
rect 87276 87502 87278 87554
rect 87330 87502 87332 87554
rect 87052 87442 87108 87454
rect 87052 87390 87054 87442
rect 87106 87390 87108 87442
rect 87052 86884 87108 87390
rect 87052 86818 87108 86828
rect 82348 85698 82404 85708
rect 82460 86546 82516 86558
rect 82460 86494 82462 86546
rect 82514 86494 82516 86546
rect 82460 86436 82516 86494
rect 85596 86548 85652 86558
rect 82124 84196 82180 84206
rect 82124 84102 82180 84140
rect 82012 83346 82068 83356
rect 82012 82738 82068 82750
rect 82012 82686 82014 82738
rect 82066 82686 82068 82738
rect 82012 82628 82068 82686
rect 82012 82562 82068 82572
rect 81452 81954 81732 81956
rect 81452 81902 81454 81954
rect 81506 81902 81732 81954
rect 81452 81900 81732 81902
rect 81452 81890 81508 81900
rect 81340 81732 81396 81742
rect 82012 81732 82068 81742
rect 80668 81678 80670 81730
rect 80722 81678 80724 81730
rect 80444 81330 80500 81340
rect 80556 81508 80612 81518
rect 80556 81394 80612 81452
rect 80556 81342 80558 81394
rect 80610 81342 80612 81394
rect 80444 81172 80500 81182
rect 80332 80836 80388 80846
rect 80332 79714 80388 80780
rect 80444 79826 80500 81116
rect 80556 81060 80612 81342
rect 80668 81284 80724 81678
rect 80668 81218 80724 81228
rect 81116 81730 81396 81732
rect 81116 81678 81342 81730
rect 81394 81678 81396 81730
rect 81116 81676 81396 81678
rect 80556 80994 80612 81004
rect 81116 80612 81172 81676
rect 81340 81666 81396 81676
rect 81788 81730 82068 81732
rect 81788 81678 82014 81730
rect 82066 81678 82068 81730
rect 81788 81676 82068 81678
rect 81276 81564 81540 81574
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81276 81498 81540 81508
rect 81452 81284 81508 81294
rect 81116 80546 81172 80556
rect 81340 81282 81508 81284
rect 81340 81230 81454 81282
rect 81506 81230 81508 81282
rect 81340 81228 81508 81230
rect 81340 80276 81396 81228
rect 81452 81218 81508 81228
rect 81676 81284 81732 81294
rect 81564 81172 81620 81182
rect 81564 81078 81620 81116
rect 81452 80948 81508 80958
rect 81452 80854 81508 80892
rect 81676 80498 81732 81228
rect 81676 80446 81678 80498
rect 81730 80446 81732 80498
rect 81676 80434 81732 80446
rect 81340 80210 81396 80220
rect 81276 79996 81540 80006
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81276 79930 81540 79940
rect 80444 79774 80446 79826
rect 80498 79774 80500 79826
rect 80444 79762 80500 79774
rect 80332 79662 80334 79714
rect 80386 79662 80388 79714
rect 80332 79650 80388 79662
rect 80668 79716 80724 79726
rect 80668 79622 80724 79660
rect 81452 79604 81508 79614
rect 81452 79510 81508 79548
rect 80444 79044 80500 79054
rect 80444 78930 80500 78988
rect 80444 78878 80446 78930
rect 80498 78878 80500 78930
rect 80444 78866 80500 78878
rect 81788 79044 81844 81676
rect 82012 81666 82068 81676
rect 82348 81284 82404 81294
rect 82348 81190 82404 81228
rect 82124 81172 82180 81182
rect 82124 81078 82180 81116
rect 82460 81170 82516 86380
rect 82572 86436 82628 86446
rect 82572 86434 82740 86436
rect 82572 86382 82574 86434
rect 82626 86382 82740 86434
rect 82572 86380 82740 86382
rect 82572 86370 82628 86380
rect 82572 85092 82628 85102
rect 82572 84998 82628 85036
rect 82684 84308 82740 86380
rect 82796 86434 82852 86446
rect 82796 86382 82798 86434
rect 82850 86382 82852 86434
rect 82796 85652 82852 86382
rect 83132 86436 83188 86446
rect 83132 86342 83188 86380
rect 84252 85874 84308 85886
rect 84252 85822 84254 85874
rect 84306 85822 84308 85874
rect 83468 85764 83524 85774
rect 84252 85764 84308 85822
rect 84812 85764 84868 85774
rect 83468 85762 83748 85764
rect 83468 85710 83470 85762
rect 83522 85710 83748 85762
rect 83468 85708 83748 85710
rect 84252 85762 84868 85764
rect 84252 85710 84814 85762
rect 84866 85710 84868 85762
rect 84252 85708 84868 85710
rect 83468 85698 83524 85708
rect 82796 85586 82852 85596
rect 83468 85092 83524 85102
rect 83020 84866 83076 84878
rect 83020 84814 83022 84866
rect 83074 84814 83076 84866
rect 83020 84308 83076 84814
rect 82684 84252 82964 84308
rect 82684 84084 82740 84094
rect 82684 82850 82740 84028
rect 82908 83636 82964 84252
rect 83020 84242 83076 84252
rect 83468 84866 83524 85036
rect 83468 84814 83470 84866
rect 83522 84814 83524 84866
rect 83020 83636 83076 83646
rect 82908 83634 83076 83636
rect 82908 83582 83022 83634
rect 83074 83582 83076 83634
rect 82908 83580 83076 83582
rect 83020 83570 83076 83580
rect 82684 82798 82686 82850
rect 82738 82798 82740 82850
rect 82684 82786 82740 82798
rect 83020 82292 83076 82302
rect 82684 81956 82740 81966
rect 82684 81862 82740 81900
rect 83020 81956 83076 82236
rect 83468 82292 83524 84814
rect 83692 83746 83748 85708
rect 84812 85092 84868 85708
rect 85596 85762 85652 86492
rect 86492 86546 86548 86558
rect 86492 86494 86494 86546
rect 86546 86494 86548 86546
rect 85596 85710 85598 85762
rect 85650 85710 85652 85762
rect 85596 85698 85652 85710
rect 86156 86434 86212 86446
rect 86156 86382 86158 86434
rect 86210 86382 86212 86434
rect 86044 85204 86100 85214
rect 86156 85204 86212 86382
rect 86492 85316 86548 86494
rect 87052 86436 87108 86446
rect 87052 86342 87108 86380
rect 87276 85988 87332 87502
rect 88396 87556 88452 87566
rect 87612 86884 87668 86894
rect 87612 86790 87668 86828
rect 87948 86658 88004 86670
rect 87948 86606 87950 86658
rect 88002 86606 88004 86658
rect 87948 86324 88004 86606
rect 88172 86546 88228 86558
rect 88172 86494 88174 86546
rect 88226 86494 88228 86546
rect 88172 86436 88228 86494
rect 88172 86370 88228 86380
rect 87948 86258 88004 86268
rect 87276 85922 87332 85932
rect 87724 85988 87780 85998
rect 87724 85894 87780 85932
rect 88396 85874 88452 87500
rect 89516 87556 89572 87566
rect 89516 87462 89572 87500
rect 90860 87556 90916 88958
rect 91644 88900 91700 88910
rect 91644 88898 91924 88900
rect 91644 88846 91646 88898
rect 91698 88846 91924 88898
rect 91644 88844 91924 88846
rect 91644 88834 91700 88844
rect 90860 87490 90916 87500
rect 88732 86548 88788 86558
rect 88732 86454 88788 86492
rect 89740 86548 89796 86558
rect 91532 86548 91588 86558
rect 88396 85822 88398 85874
rect 88450 85822 88452 85874
rect 88396 85810 88452 85822
rect 89180 86436 89236 86446
rect 86492 85250 86548 85260
rect 88060 85764 88116 85774
rect 86044 85202 86212 85204
rect 86044 85150 86046 85202
rect 86098 85150 86212 85202
rect 86044 85148 86212 85150
rect 87500 85204 87556 85214
rect 86044 85138 86100 85148
rect 85372 85092 85428 85102
rect 84812 85090 85428 85092
rect 84812 85038 85374 85090
rect 85426 85038 85428 85090
rect 84812 85036 85428 85038
rect 84924 84420 84980 84430
rect 84924 84326 84980 84364
rect 85036 84306 85092 84318
rect 85036 84254 85038 84306
rect 85090 84254 85092 84306
rect 83692 83694 83694 83746
rect 83746 83694 83748 83746
rect 83692 83682 83748 83694
rect 84252 84194 84308 84206
rect 84252 84142 84254 84194
rect 84306 84142 84308 84194
rect 83580 83412 83636 83422
rect 83580 83318 83636 83356
rect 83692 83300 83748 83310
rect 83692 83298 83860 83300
rect 83692 83246 83694 83298
rect 83746 83246 83860 83298
rect 83692 83244 83860 83246
rect 83692 83234 83748 83244
rect 83468 82226 83524 82236
rect 83020 81954 83300 81956
rect 83020 81902 83022 81954
rect 83074 81902 83300 81954
rect 83020 81900 83300 81902
rect 83020 81890 83076 81900
rect 83244 81844 83300 81900
rect 83580 81844 83636 81854
rect 83244 81842 83636 81844
rect 83244 81790 83582 81842
rect 83634 81790 83636 81842
rect 83244 81788 83636 81790
rect 82908 81730 82964 81742
rect 82908 81678 82910 81730
rect 82962 81678 82964 81730
rect 82908 81620 82964 81678
rect 82908 81554 82964 81564
rect 83132 81282 83188 81294
rect 83132 81230 83134 81282
rect 83186 81230 83188 81282
rect 82460 81118 82462 81170
rect 82514 81118 82516 81170
rect 82460 81060 82516 81118
rect 82460 80994 82516 81004
rect 82908 81170 82964 81182
rect 82908 81118 82910 81170
rect 82962 81118 82964 81170
rect 82908 80836 82964 81118
rect 82908 80770 82964 80780
rect 81276 78428 81540 78438
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81276 78362 81540 78372
rect 80332 78036 80388 78046
rect 80220 78034 80388 78036
rect 80220 77982 80334 78034
rect 80386 77982 80388 78034
rect 80220 77980 80388 77982
rect 80220 76690 80276 77980
rect 80332 77970 80388 77980
rect 81452 78034 81508 78046
rect 81452 77982 81454 78034
rect 81506 77982 81508 78034
rect 81340 77924 81396 77934
rect 80780 77364 80836 77374
rect 80444 77252 80500 77262
rect 80444 77158 80500 77196
rect 80780 77250 80836 77308
rect 80780 77198 80782 77250
rect 80834 77198 80836 77250
rect 80220 76638 80222 76690
rect 80274 76638 80276 76690
rect 80220 76626 80276 76638
rect 80780 76692 80836 77198
rect 81340 77140 81396 77868
rect 81452 77364 81508 77982
rect 81788 77364 81844 78988
rect 82012 80724 82068 80734
rect 82012 78818 82068 80668
rect 82908 80388 82964 80398
rect 82908 80294 82964 80332
rect 83020 80276 83076 80286
rect 82236 80164 82292 80174
rect 82236 80070 82292 80108
rect 82572 80162 82628 80174
rect 82572 80110 82574 80162
rect 82626 80110 82628 80162
rect 82124 79716 82180 79726
rect 82124 79622 82180 79660
rect 82572 78988 82628 80110
rect 82012 78766 82014 78818
rect 82066 78766 82068 78818
rect 82012 78754 82068 78766
rect 82348 78932 82628 78988
rect 82796 80162 82852 80174
rect 82796 80110 82798 80162
rect 82850 80110 82852 80162
rect 82124 77924 82180 77934
rect 82124 77830 82180 77868
rect 82236 77364 82292 77374
rect 81452 77362 82292 77364
rect 81452 77310 82238 77362
rect 82290 77310 82292 77362
rect 81452 77308 82292 77310
rect 82236 77298 82292 77308
rect 81452 77140 81508 77150
rect 81340 77138 81508 77140
rect 81340 77086 81454 77138
rect 81506 77086 81508 77138
rect 81340 77084 81508 77086
rect 81452 77074 81508 77084
rect 81788 77140 81844 77150
rect 82348 77140 82404 78932
rect 82796 78820 82852 80110
rect 82796 78754 82852 78764
rect 83020 78818 83076 80220
rect 83132 79492 83188 81230
rect 83244 81282 83300 81788
rect 83580 81778 83636 81788
rect 83692 81732 83748 81742
rect 83692 81638 83748 81676
rect 83244 81230 83246 81282
rect 83298 81230 83300 81282
rect 83244 81218 83300 81230
rect 83692 81060 83748 81070
rect 83580 80612 83636 80622
rect 83580 80518 83636 80556
rect 83580 80276 83636 80286
rect 83468 80220 83580 80276
rect 83132 79426 83188 79436
rect 83244 80164 83300 80174
rect 83020 78766 83022 78818
rect 83074 78766 83076 78818
rect 83020 78754 83076 78766
rect 83132 79268 83188 79278
rect 83020 77140 83076 77150
rect 81788 77138 82404 77140
rect 81788 77086 81790 77138
rect 81842 77086 82404 77138
rect 81788 77084 82404 77086
rect 82908 77084 83020 77140
rect 81788 77074 81844 77084
rect 81676 77026 81732 77038
rect 81676 76974 81678 77026
rect 81730 76974 81732 77026
rect 81276 76860 81540 76870
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81276 76794 81540 76804
rect 80780 76626 80836 76636
rect 81452 76578 81508 76590
rect 81452 76526 81454 76578
rect 81506 76526 81508 76578
rect 80556 76468 80612 76478
rect 80556 76354 80612 76412
rect 80556 76302 80558 76354
rect 80610 76302 80612 76354
rect 79772 75796 79828 75806
rect 79772 75702 79828 75740
rect 80556 75572 80612 76302
rect 81228 76466 81284 76478
rect 81228 76414 81230 76466
rect 81282 76414 81284 76466
rect 81228 75796 81284 76414
rect 81228 75730 81284 75740
rect 81452 75684 81508 76526
rect 81564 76468 81620 76478
rect 81676 76468 81732 76974
rect 82236 76580 82292 76590
rect 81564 76466 81732 76468
rect 81564 76414 81566 76466
rect 81618 76414 81732 76466
rect 81564 76412 81732 76414
rect 81900 76578 82292 76580
rect 81900 76526 82238 76578
rect 82290 76526 82292 76578
rect 81900 76524 82292 76526
rect 81564 76244 81620 76412
rect 81564 76178 81620 76188
rect 81900 75794 81956 76524
rect 82236 76514 82292 76524
rect 82796 76580 82852 76590
rect 82908 76580 82964 77084
rect 83020 77008 83076 77084
rect 83132 77138 83188 79212
rect 83132 77086 83134 77138
rect 83186 77086 83188 77138
rect 82852 76524 82964 76580
rect 82348 76468 82404 76478
rect 82348 76374 82404 76412
rect 82236 76244 82292 76254
rect 82236 76150 82292 76188
rect 81900 75742 81902 75794
rect 81954 75742 81956 75794
rect 81900 75730 81956 75742
rect 81452 75618 81508 75628
rect 82348 75684 82404 75694
rect 82348 75590 82404 75628
rect 82684 75684 82740 75694
rect 82796 75684 82852 76524
rect 83132 75684 83188 77086
rect 83244 78594 83300 80108
rect 83468 79268 83524 80220
rect 83580 80182 83636 80220
rect 83692 80274 83748 81004
rect 83692 80222 83694 80274
rect 83746 80222 83748 80274
rect 83468 79202 83524 79212
rect 83580 79604 83636 79614
rect 83580 78932 83636 79548
rect 83356 78708 83412 78718
rect 83356 78614 83412 78652
rect 83244 78542 83246 78594
rect 83298 78542 83300 78594
rect 83244 75796 83300 78542
rect 83356 77028 83412 77038
rect 83356 76934 83412 76972
rect 83580 76466 83636 78876
rect 83692 78708 83748 80222
rect 83804 78818 83860 83244
rect 83916 82740 83972 82750
rect 83916 81954 83972 82684
rect 83916 81902 83918 81954
rect 83970 81902 83972 81954
rect 83916 81890 83972 81902
rect 84140 82292 84196 82302
rect 84140 81058 84196 82236
rect 84252 81620 84308 84142
rect 84924 84084 84980 84094
rect 84924 83990 84980 84028
rect 84364 83300 84420 83310
rect 84364 83298 84532 83300
rect 84364 83246 84366 83298
rect 84418 83246 84532 83298
rect 84364 83244 84532 83246
rect 84364 83234 84420 83244
rect 84252 81554 84308 81564
rect 84364 81730 84420 81742
rect 84364 81678 84366 81730
rect 84418 81678 84420 81730
rect 84140 81006 84142 81058
rect 84194 81006 84196 81058
rect 84140 80724 84196 81006
rect 84364 81060 84420 81678
rect 84364 80994 84420 81004
rect 84140 80658 84196 80668
rect 84252 80388 84308 80398
rect 84252 80294 84308 80332
rect 84476 80276 84532 83244
rect 85036 82740 85092 84254
rect 85260 83300 85316 83310
rect 85036 82674 85092 82684
rect 85148 83298 85316 83300
rect 85148 83246 85262 83298
rect 85314 83246 85316 83298
rect 85148 83244 85316 83246
rect 84812 82626 84868 82638
rect 84812 82574 84814 82626
rect 84866 82574 84868 82626
rect 84812 81732 84868 82574
rect 84588 81060 84644 81070
rect 84588 80966 84644 81004
rect 84812 80836 84868 81676
rect 85148 80948 85204 83244
rect 85260 83234 85316 83244
rect 85260 82628 85316 82638
rect 85372 82628 85428 85036
rect 85596 84194 85652 84206
rect 85596 84142 85598 84194
rect 85650 84142 85652 84194
rect 85596 83748 85652 84142
rect 85596 83682 85652 83692
rect 87388 83748 87444 83758
rect 85316 82572 85428 82628
rect 85708 83298 85764 83310
rect 85708 83246 85710 83298
rect 85762 83246 85764 83298
rect 85260 82534 85316 82572
rect 85708 82514 85764 83246
rect 85708 82462 85710 82514
rect 85762 82462 85764 82514
rect 85708 82450 85764 82462
rect 85820 82628 85876 82638
rect 86156 82628 86212 82638
rect 85820 82626 86212 82628
rect 85820 82574 85822 82626
rect 85874 82574 86158 82626
rect 86210 82574 86212 82626
rect 85820 82572 86212 82574
rect 85260 81620 85316 81630
rect 85260 81282 85316 81564
rect 85260 81230 85262 81282
rect 85314 81230 85316 81282
rect 85260 81218 85316 81230
rect 85708 81172 85764 81182
rect 85820 81172 85876 82572
rect 86156 82562 86212 82572
rect 86604 82628 86660 82638
rect 86604 82534 86660 82572
rect 86716 82516 86772 82526
rect 86716 82514 86884 82516
rect 86716 82462 86718 82514
rect 86770 82462 86884 82514
rect 86716 82460 86884 82462
rect 86716 82450 86772 82460
rect 86716 81954 86772 81966
rect 86716 81902 86718 81954
rect 86770 81902 86772 81954
rect 86268 81284 86324 81294
rect 86268 81282 86660 81284
rect 86268 81230 86270 81282
rect 86322 81230 86660 81282
rect 86268 81228 86660 81230
rect 86268 81218 86324 81228
rect 86044 81172 86100 81182
rect 85708 81170 85876 81172
rect 85708 81118 85710 81170
rect 85762 81118 85876 81170
rect 85708 81116 85876 81118
rect 85708 81106 85764 81116
rect 85148 80892 85652 80948
rect 84812 80780 85316 80836
rect 84476 80210 84532 80220
rect 84700 80276 84756 80286
rect 84364 80162 84420 80174
rect 84364 80110 84366 80162
rect 84418 80110 84420 80162
rect 84364 79604 84420 80110
rect 84364 79538 84420 79548
rect 84588 80162 84644 80174
rect 84588 80110 84590 80162
rect 84642 80110 84644 80162
rect 84252 79492 84308 79502
rect 84252 79398 84308 79436
rect 84476 79378 84532 79390
rect 84476 79326 84478 79378
rect 84530 79326 84532 79378
rect 84476 78988 84532 79326
rect 83804 78766 83806 78818
rect 83858 78766 83860 78818
rect 83804 78754 83860 78766
rect 84028 78932 84532 78988
rect 83692 78642 83748 78652
rect 84028 78706 84084 78932
rect 84252 78820 84308 78830
rect 84028 78654 84030 78706
rect 84082 78654 84084 78706
rect 84028 77252 84084 78654
rect 84140 78708 84196 78718
rect 84140 78614 84196 78652
rect 84252 77922 84308 78764
rect 84588 78148 84644 80110
rect 84700 79826 84756 80220
rect 85148 80164 85204 80174
rect 84700 79774 84702 79826
rect 84754 79774 84756 79826
rect 84700 79762 84756 79774
rect 85036 80162 85204 80164
rect 85036 80110 85150 80162
rect 85202 80110 85204 80162
rect 85036 80108 85204 80110
rect 85036 79378 85092 80108
rect 85148 80098 85204 80108
rect 85260 79714 85316 80780
rect 85596 80498 85652 80892
rect 85596 80446 85598 80498
rect 85650 80446 85652 80498
rect 85260 79662 85262 79714
rect 85314 79662 85316 79714
rect 85260 79650 85316 79662
rect 85372 80388 85428 80398
rect 85036 79326 85038 79378
rect 85090 79326 85092 79378
rect 85036 79314 85092 79326
rect 85260 79492 85316 79502
rect 85260 78930 85316 79436
rect 85260 78878 85262 78930
rect 85314 78878 85316 78930
rect 85260 78866 85316 78878
rect 84588 78082 84644 78092
rect 84252 77870 84254 77922
rect 84306 77870 84308 77922
rect 84252 77858 84308 77870
rect 84700 77922 84756 77934
rect 84700 77870 84702 77922
rect 84754 77870 84756 77922
rect 83916 77196 84084 77252
rect 84364 77364 84420 77374
rect 84364 77250 84420 77308
rect 84364 77198 84366 77250
rect 84418 77198 84420 77250
rect 83916 76804 83972 77196
rect 84364 77186 84420 77198
rect 84700 77140 84756 77870
rect 85260 77362 85316 77374
rect 85260 77310 85262 77362
rect 85314 77310 85316 77362
rect 85260 77252 85316 77310
rect 85260 77186 85316 77196
rect 84700 77074 84756 77084
rect 84028 77028 84084 77038
rect 84252 77028 84308 77038
rect 84028 77026 84196 77028
rect 84028 76974 84030 77026
rect 84082 76974 84196 77026
rect 84028 76972 84196 76974
rect 84028 76962 84084 76972
rect 83916 76748 84084 76804
rect 83580 76414 83582 76466
rect 83634 76414 83636 76466
rect 83580 76402 83636 76414
rect 83244 75740 83412 75796
rect 82684 75682 82796 75684
rect 82684 75630 82686 75682
rect 82738 75630 82796 75682
rect 82684 75628 82796 75630
rect 80556 75506 80612 75516
rect 82236 75460 82292 75470
rect 81276 75292 81540 75302
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81276 75226 81540 75236
rect 81788 74898 81844 74910
rect 81788 74846 81790 74898
rect 81842 74846 81844 74898
rect 81340 74788 81396 74798
rect 81788 74788 81844 74846
rect 78764 73892 78932 73948
rect 78764 73444 78820 73454
rect 78764 73350 78820 73388
rect 78652 69682 78708 69692
rect 78204 69410 78260 69422
rect 78204 69358 78206 69410
rect 78258 69358 78260 69410
rect 77980 69300 78036 69310
rect 77756 69298 78036 69300
rect 77756 69246 77982 69298
rect 78034 69246 78036 69298
rect 77756 69244 78036 69246
rect 77420 69206 77476 69244
rect 77196 68798 77198 68850
rect 77250 68798 77252 68850
rect 77196 68786 77252 68798
rect 77756 68626 77812 68638
rect 77756 68574 77758 68626
rect 77810 68574 77812 68626
rect 77084 68012 77252 68068
rect 77196 67956 77252 68012
rect 77532 67956 77588 67966
rect 77196 67954 77588 67956
rect 77196 67902 77534 67954
rect 77586 67902 77588 67954
rect 77196 67900 77588 67902
rect 77420 67732 77476 67742
rect 77084 67170 77140 67182
rect 77084 67118 77086 67170
rect 77138 67118 77140 67170
rect 76748 67058 76804 67070
rect 76748 67006 76750 67058
rect 76802 67006 76804 67058
rect 76748 66948 76804 67006
rect 77084 67060 77140 67118
rect 77084 66994 77140 67004
rect 76748 66882 76804 66892
rect 77420 66500 77476 67676
rect 77532 67060 77588 67900
rect 77644 67060 77700 67070
rect 77532 67058 77700 67060
rect 77532 67006 77646 67058
rect 77698 67006 77700 67058
rect 77532 67004 77700 67006
rect 77420 66274 77476 66444
rect 77420 66222 77422 66274
rect 77474 66222 77476 66274
rect 77196 65490 77252 65502
rect 77196 65438 77198 65490
rect 77250 65438 77252 65490
rect 77196 64708 77252 65438
rect 77196 64652 77364 64708
rect 76524 63410 76580 63420
rect 76860 64484 76916 64494
rect 76412 63086 76414 63138
rect 76466 63086 76468 63138
rect 76412 63074 76468 63086
rect 76300 61842 76356 61852
rect 76412 62914 76468 62926
rect 76412 62862 76414 62914
rect 76466 62862 76468 62914
rect 75852 61518 75854 61570
rect 75906 61518 75908 61570
rect 75852 61506 75908 61518
rect 75964 61346 76020 61358
rect 75964 61294 75966 61346
rect 76018 61294 76020 61346
rect 75852 60116 75908 60126
rect 75852 60022 75908 60060
rect 75852 59220 75908 59230
rect 75740 59218 75908 59220
rect 75740 59166 75854 59218
rect 75906 59166 75908 59218
rect 75740 59164 75908 59166
rect 75852 59108 75908 59164
rect 75852 59042 75908 59052
rect 75628 58436 75684 58446
rect 75628 58342 75684 58380
rect 75852 58212 75908 58222
rect 75516 58034 75572 58044
rect 75740 58210 75908 58212
rect 75740 58158 75854 58210
rect 75906 58158 75908 58210
rect 75740 58156 75908 58158
rect 75404 57698 75460 57708
rect 75740 57652 75796 58156
rect 75852 58146 75908 58156
rect 75852 57764 75908 57774
rect 75852 57670 75908 57708
rect 75628 57650 75796 57652
rect 75628 57598 75742 57650
rect 75794 57598 75796 57650
rect 75628 57596 75796 57598
rect 75292 57092 75348 57102
rect 75292 56868 75348 57036
rect 75628 56868 75684 57596
rect 75740 57586 75796 57596
rect 75964 56980 76020 61294
rect 76300 61346 76356 61358
rect 76300 61294 76302 61346
rect 76354 61294 76356 61346
rect 76300 61236 76356 61294
rect 76300 61170 76356 61180
rect 76412 60116 76468 62862
rect 76300 60060 76468 60116
rect 76524 62916 76580 62926
rect 76524 60116 76580 62860
rect 76860 62580 76916 64428
rect 77196 64482 77252 64494
rect 77196 64430 77198 64482
rect 77250 64430 77252 64482
rect 77196 64372 77252 64430
rect 76860 62514 76916 62524
rect 76972 64316 77252 64372
rect 76972 61460 77028 64316
rect 77308 64260 77364 64652
rect 77084 64204 77364 64260
rect 77084 64036 77140 64204
rect 77084 63922 77140 63980
rect 77084 63870 77086 63922
rect 77138 63870 77140 63922
rect 77084 63858 77140 63870
rect 77196 63924 77252 63934
rect 77196 62188 77252 63868
rect 77308 63252 77364 63262
rect 77308 63158 77364 63196
rect 77196 62132 77364 62188
rect 77308 61572 77364 62132
rect 77308 61478 77364 61516
rect 76748 60676 76804 60686
rect 76748 60582 76804 60620
rect 76972 60228 77028 61404
rect 77420 61348 77476 66222
rect 77644 66276 77700 67004
rect 77644 66210 77700 66220
rect 77756 66164 77812 68574
rect 77980 68628 78036 69244
rect 78204 69300 78260 69358
rect 78204 69234 78260 69244
rect 78540 69188 78596 69198
rect 78540 69094 78596 69132
rect 78876 68852 78932 73892
rect 79212 73892 79492 73948
rect 81116 74786 81844 74788
rect 81116 74734 81342 74786
rect 81394 74734 81844 74786
rect 81116 74732 81844 74734
rect 78988 73108 79044 73118
rect 78988 73014 79044 73052
rect 78988 72434 79044 72446
rect 78988 72382 78990 72434
rect 79042 72382 79044 72434
rect 78988 72212 79044 72382
rect 78988 72146 79044 72156
rect 79100 72324 79156 72334
rect 79100 69412 79156 72268
rect 79100 69318 79156 69356
rect 79212 69076 79268 73892
rect 79324 73556 79380 73566
rect 79324 73462 79380 73500
rect 79996 73218 80052 73230
rect 79996 73166 79998 73218
rect 80050 73166 80052 73218
rect 79996 73108 80052 73166
rect 79996 71652 80052 73052
rect 79996 71586 80052 71596
rect 80332 72212 80388 72222
rect 80332 71092 80388 72156
rect 81116 72212 81172 74732
rect 81340 74722 81396 74732
rect 82236 74228 82292 75404
rect 82572 75460 82628 75470
rect 82572 75366 82628 75404
rect 82572 74786 82628 74798
rect 82572 74734 82574 74786
rect 82626 74734 82628 74786
rect 82572 74338 82628 74734
rect 82572 74286 82574 74338
rect 82626 74286 82628 74338
rect 82572 74274 82628 74286
rect 82236 74096 82292 74172
rect 82684 74226 82740 75628
rect 82796 75552 82852 75628
rect 83020 75628 83188 75684
rect 83020 74564 83076 75628
rect 83244 75572 83300 75582
rect 83020 74498 83076 74508
rect 83132 75458 83188 75470
rect 83132 75406 83134 75458
rect 83186 75406 83188 75458
rect 82908 74340 82964 74350
rect 82908 74338 83076 74340
rect 82908 74286 82910 74338
rect 82962 74286 83076 74338
rect 82908 74284 83076 74286
rect 82908 74274 82964 74284
rect 82684 74174 82686 74226
rect 82738 74174 82740 74226
rect 82684 74162 82740 74174
rect 82796 74228 82852 74238
rect 81276 73724 81540 73734
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81276 73658 81540 73668
rect 81788 73444 81844 73454
rect 81788 73442 82180 73444
rect 81788 73390 81790 73442
rect 81842 73390 82180 73442
rect 81788 73388 82180 73390
rect 81788 73378 81844 73388
rect 81564 73332 81620 73342
rect 81564 73330 81732 73332
rect 81564 73278 81566 73330
rect 81618 73278 81732 73330
rect 81564 73276 81732 73278
rect 81564 73266 81620 73276
rect 81116 71764 81172 72156
rect 81276 72156 81540 72166
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81276 72090 81540 72100
rect 81340 71764 81396 71774
rect 81116 71762 81396 71764
rect 81116 71710 81342 71762
rect 81394 71710 81396 71762
rect 81116 71708 81396 71710
rect 81340 71698 81396 71708
rect 80556 71652 80612 71662
rect 80556 71558 80612 71596
rect 81564 71652 81620 71662
rect 80780 71092 80836 71102
rect 80332 71090 81172 71092
rect 80332 71038 80334 71090
rect 80386 71038 80782 71090
rect 80834 71038 81172 71090
rect 80332 71036 81172 71038
rect 80332 71026 80388 71036
rect 80780 71026 80836 71036
rect 81116 70420 81172 71036
rect 81564 70868 81620 71596
rect 81676 71204 81732 73276
rect 82124 71874 82180 73388
rect 82124 71822 82126 71874
rect 82178 71822 82180 71874
rect 82124 71810 82180 71822
rect 82012 71204 82068 71214
rect 81676 71202 82068 71204
rect 81676 71150 82014 71202
rect 82066 71150 82068 71202
rect 81676 71148 82068 71150
rect 82012 71138 82068 71148
rect 82348 71204 82404 71214
rect 82348 71110 82404 71148
rect 82796 70868 82852 74172
rect 83020 74114 83076 74284
rect 83020 74062 83022 74114
rect 83074 74062 83076 74114
rect 83020 74050 83076 74062
rect 83132 73892 83188 75406
rect 83244 74116 83300 75516
rect 83356 75458 83412 75740
rect 83468 75684 83524 75694
rect 83468 75590 83524 75628
rect 83356 75406 83358 75458
rect 83410 75406 83412 75458
rect 83356 75236 83412 75406
rect 84028 75460 84084 76748
rect 84140 76580 84196 76972
rect 84252 76934 84308 76972
rect 85372 76916 85428 80332
rect 85596 80388 85652 80446
rect 85596 80322 85652 80332
rect 85708 80610 85764 80622
rect 85708 80558 85710 80610
rect 85762 80558 85764 80610
rect 85596 80052 85652 80062
rect 85484 79604 85540 79614
rect 85484 77922 85540 79548
rect 85596 79602 85652 79996
rect 85596 79550 85598 79602
rect 85650 79550 85652 79602
rect 85596 79538 85652 79550
rect 85484 77870 85486 77922
rect 85538 77870 85540 77922
rect 85484 77858 85540 77870
rect 85708 78818 85764 80558
rect 85820 80052 85876 81116
rect 85820 79986 85876 79996
rect 85932 81170 86100 81172
rect 85932 81118 86046 81170
rect 86098 81118 86100 81170
rect 85932 81116 86100 81118
rect 85708 78766 85710 78818
rect 85762 78766 85764 78818
rect 85372 76850 85428 76860
rect 85596 77364 85652 77374
rect 84252 76580 84308 76590
rect 84140 76578 84308 76580
rect 84140 76526 84254 76578
rect 84306 76526 84308 76578
rect 84140 76524 84308 76526
rect 84252 76514 84308 76524
rect 84028 75394 84084 75404
rect 84252 76356 84308 76366
rect 84252 75684 84308 76300
rect 85372 76356 85428 76366
rect 84252 75570 84308 75628
rect 84252 75518 84254 75570
rect 84306 75518 84308 75570
rect 83356 75180 83860 75236
rect 83580 74564 83636 74574
rect 83356 74116 83412 74126
rect 83244 74114 83412 74116
rect 83244 74062 83358 74114
rect 83410 74062 83412 74114
rect 83244 74060 83412 74062
rect 83356 74050 83412 74060
rect 83244 73892 83300 73902
rect 83132 73890 83300 73892
rect 83132 73838 83246 73890
rect 83298 73838 83300 73890
rect 83132 73836 83300 73838
rect 83244 73826 83300 73836
rect 83244 73442 83300 73454
rect 83244 73390 83246 73442
rect 83298 73390 83300 73442
rect 83020 73330 83076 73342
rect 83020 73278 83022 73330
rect 83074 73278 83076 73330
rect 83020 71876 83076 73278
rect 83020 71810 83076 71820
rect 83020 70978 83076 70990
rect 83020 70926 83022 70978
rect 83074 70926 83076 70978
rect 82908 70868 82964 70878
rect 81564 70812 81732 70868
rect 81452 70756 81508 70794
rect 81452 70690 81508 70700
rect 81276 70588 81540 70598
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81276 70522 81540 70532
rect 81228 70420 81284 70430
rect 81116 70418 81284 70420
rect 81116 70366 81230 70418
rect 81282 70366 81284 70418
rect 81116 70364 81284 70366
rect 81228 70354 81284 70364
rect 80444 70082 80500 70094
rect 80444 70030 80446 70082
rect 80498 70030 80500 70082
rect 79996 69300 80052 69310
rect 78764 68796 78932 68852
rect 78988 69020 79268 69076
rect 79548 69186 79604 69198
rect 79548 69134 79550 69186
rect 79602 69134 79604 69186
rect 78092 68740 78148 68750
rect 78092 68646 78148 68684
rect 77980 68068 78036 68572
rect 77980 68002 78036 68012
rect 78652 68514 78708 68526
rect 78652 68462 78654 68514
rect 78706 68462 78708 68514
rect 77644 66050 77700 66062
rect 77644 65998 77646 66050
rect 77698 65998 77700 66050
rect 77532 65940 77588 65950
rect 77644 65940 77700 65998
rect 77588 65884 77700 65940
rect 77532 65874 77588 65884
rect 77756 65828 77812 66108
rect 78428 66946 78484 66958
rect 78428 66894 78430 66946
rect 78482 66894 78484 66946
rect 77644 65772 77812 65828
rect 77868 66052 77924 66062
rect 77644 64146 77700 65772
rect 77756 65604 77812 65614
rect 77868 65604 77924 65996
rect 77756 65602 77924 65604
rect 77756 65550 77758 65602
rect 77810 65550 77924 65602
rect 77756 65548 77924 65550
rect 77756 65538 77812 65548
rect 78092 65492 78148 65502
rect 78428 65492 78484 66894
rect 78652 66388 78708 68462
rect 78652 66322 78708 66332
rect 78540 66276 78596 66286
rect 78540 66182 78596 66220
rect 78092 65490 78260 65492
rect 78092 65438 78094 65490
rect 78146 65438 78260 65490
rect 78092 65436 78260 65438
rect 78092 65426 78148 65436
rect 78092 65044 78148 65054
rect 77868 64484 77924 64494
rect 77868 64390 77924 64428
rect 77644 64094 77646 64146
rect 77698 64094 77700 64146
rect 77644 64082 77700 64094
rect 77756 64148 77812 64158
rect 78092 64148 78148 64988
rect 78204 64596 78260 65436
rect 78428 65426 78484 65436
rect 78540 65828 78596 65838
rect 78540 65380 78596 65772
rect 78316 64596 78372 64606
rect 78204 64594 78316 64596
rect 78204 64542 78206 64594
rect 78258 64542 78316 64594
rect 78204 64540 78316 64542
rect 78204 64530 78260 64540
rect 78204 64148 78260 64158
rect 78092 64146 78260 64148
rect 78092 64094 78206 64146
rect 78258 64094 78260 64146
rect 78092 64092 78260 64094
rect 77756 64034 77812 64092
rect 78204 64082 78260 64092
rect 77756 63982 77758 64034
rect 77810 63982 77812 64034
rect 77756 63364 77812 63982
rect 77980 63924 78036 63934
rect 77980 63830 78036 63868
rect 77756 63298 77812 63308
rect 77868 63700 77924 63710
rect 77756 63140 77812 63150
rect 77420 61282 77476 61292
rect 77532 63138 77812 63140
rect 77532 63086 77758 63138
rect 77810 63086 77812 63138
rect 77532 63084 77812 63086
rect 77532 62466 77588 63084
rect 77756 63074 77812 63084
rect 77532 62414 77534 62466
rect 77586 62414 77588 62466
rect 77532 60452 77588 62414
rect 77868 62188 77924 63644
rect 78316 62580 78372 64540
rect 78428 64036 78484 64046
rect 78540 64036 78596 65324
rect 78428 64034 78596 64036
rect 78428 63982 78430 64034
rect 78482 63982 78596 64034
rect 78428 63980 78596 63982
rect 78428 63970 78484 63980
rect 78764 63812 78820 68796
rect 78876 65490 78932 65502
rect 78876 65438 78878 65490
rect 78930 65438 78932 65490
rect 78876 64596 78932 65438
rect 78988 64932 79044 69020
rect 79548 68964 79604 69134
rect 79996 69188 80052 69244
rect 80444 69188 80500 70030
rect 81228 69524 81284 69534
rect 81228 69430 81284 69468
rect 79996 69186 80500 69188
rect 79996 69134 79998 69186
rect 80050 69134 80500 69186
rect 79996 69132 80500 69134
rect 79996 69122 80052 69132
rect 79100 68908 79604 68964
rect 79100 68740 79156 68908
rect 79100 68626 79156 68684
rect 79100 68574 79102 68626
rect 79154 68574 79156 68626
rect 79100 67620 79156 68574
rect 79100 67554 79156 67564
rect 79212 68738 79268 68750
rect 79212 68686 79214 68738
rect 79266 68686 79268 68738
rect 79212 66948 79268 68686
rect 79996 68740 80052 68750
rect 79996 68738 80164 68740
rect 79996 68686 79998 68738
rect 80050 68686 80164 68738
rect 79996 68684 80164 68686
rect 79996 68674 80052 68684
rect 79436 68628 79492 68638
rect 79884 68628 79940 68638
rect 79436 68626 79940 68628
rect 79436 68574 79438 68626
rect 79490 68574 79886 68626
rect 79938 68574 79940 68626
rect 79436 68572 79940 68574
rect 79436 68562 79492 68572
rect 79212 66882 79268 66892
rect 79324 68404 79380 68414
rect 79100 66612 79156 66622
rect 79100 65716 79156 66556
rect 79324 66386 79380 68348
rect 79324 66334 79326 66386
rect 79378 66334 79380 66386
rect 79324 66322 79380 66334
rect 79100 65584 79156 65660
rect 79772 65714 79828 68572
rect 79884 68562 79940 68572
rect 79996 68404 80052 68414
rect 79996 68310 80052 68348
rect 80108 67172 80164 68684
rect 80108 67106 80164 67116
rect 80220 66948 80276 69132
rect 81276 69020 81540 69030
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81276 68954 81540 68964
rect 81276 67452 81540 67462
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81276 67386 81540 67396
rect 81228 67172 81284 67182
rect 81228 67078 81284 67116
rect 81452 67170 81508 67182
rect 81452 67118 81454 67170
rect 81506 67118 81508 67170
rect 79772 65662 79774 65714
rect 79826 65662 79828 65714
rect 79772 65650 79828 65662
rect 79884 66892 80276 66948
rect 80556 66948 80612 66958
rect 79660 65604 79716 65614
rect 79660 65510 79716 65548
rect 79884 65492 79940 66892
rect 80556 66854 80612 66892
rect 80668 66836 80724 66846
rect 80668 65940 80724 66780
rect 79772 65436 79940 65492
rect 79996 65492 80052 65502
rect 79660 65156 79716 65166
rect 78988 64820 79044 64876
rect 79436 65044 79492 65054
rect 78988 64764 79156 64820
rect 78988 64596 79044 64606
rect 78876 64540 78988 64596
rect 78988 64502 79044 64540
rect 79100 64148 79156 64764
rect 79324 64482 79380 64494
rect 79324 64430 79326 64482
rect 79378 64430 79380 64482
rect 79324 64372 79380 64430
rect 79100 64082 79156 64092
rect 79212 64316 79324 64372
rect 78764 63746 78820 63756
rect 78988 63922 79044 63934
rect 78988 63870 78990 63922
rect 79042 63870 79044 63922
rect 78540 63140 78596 63150
rect 78428 62580 78484 62590
rect 78316 62578 78484 62580
rect 78316 62526 78430 62578
rect 78482 62526 78484 62578
rect 78316 62524 78484 62526
rect 78428 62514 78484 62524
rect 78092 62354 78148 62366
rect 78092 62302 78094 62354
rect 78146 62302 78148 62354
rect 77868 62132 78036 62188
rect 77980 61460 78036 62132
rect 77980 61394 78036 61404
rect 78092 62132 78148 62302
rect 78540 62188 78596 63084
rect 78764 63028 78820 63038
rect 78764 62934 78820 62972
rect 77868 61346 77924 61358
rect 77868 61294 77870 61346
rect 77922 61294 77924 61346
rect 77868 61012 77924 61294
rect 77868 60946 77924 60956
rect 77532 60386 77588 60396
rect 76972 60162 77028 60172
rect 77644 60228 77700 60238
rect 76188 58996 76244 59006
rect 76076 58548 76132 58558
rect 76076 58434 76132 58492
rect 76076 58382 76078 58434
rect 76130 58382 76132 58434
rect 76076 58370 76132 58382
rect 76188 57874 76244 58940
rect 76188 57822 76190 57874
rect 76242 57822 76244 57874
rect 76188 57810 76244 57822
rect 76300 56980 76356 60060
rect 76524 60050 76580 60060
rect 76412 59892 76468 59902
rect 76412 59798 76468 59836
rect 77644 59890 77700 60172
rect 77644 59838 77646 59890
rect 77698 59838 77700 59890
rect 77644 59826 77700 59838
rect 78092 60004 78148 62076
rect 77308 59780 77364 59790
rect 77308 59686 77364 59724
rect 77532 59668 77588 59678
rect 76972 59330 77028 59342
rect 76972 59278 76974 59330
rect 77026 59278 77028 59330
rect 76972 58996 77028 59278
rect 76972 58930 77028 58940
rect 77084 58324 77140 58334
rect 76524 58212 76580 58222
rect 76524 58118 76580 58156
rect 76972 57876 77028 57886
rect 76860 57764 76916 57774
rect 76860 57670 76916 57708
rect 76972 57762 77028 57820
rect 76972 57710 76974 57762
rect 77026 57710 77028 57762
rect 76972 57698 77028 57710
rect 77084 57764 77140 58268
rect 77308 58322 77364 58334
rect 77308 58270 77310 58322
rect 77362 58270 77364 58322
rect 77084 57698 77140 57708
rect 77196 58212 77252 58222
rect 76524 57652 76580 57662
rect 76412 56980 76468 56990
rect 75964 56924 76132 56980
rect 75292 56812 76020 56868
rect 75292 56754 75348 56812
rect 75292 56702 75294 56754
rect 75346 56702 75348 56754
rect 75292 56690 75348 56702
rect 75964 56754 76020 56812
rect 75964 56702 75966 56754
rect 76018 56702 76020 56754
rect 75964 56690 76020 56702
rect 75404 56644 75460 56654
rect 75404 56306 75460 56588
rect 75404 56254 75406 56306
rect 75458 56254 75460 56306
rect 75404 56242 75460 56254
rect 75852 56642 75908 56654
rect 75852 56590 75854 56642
rect 75906 56590 75908 56642
rect 75852 56196 75908 56590
rect 75740 56084 75796 56094
rect 75740 55990 75796 56028
rect 75852 55524 75908 56140
rect 75852 55458 75908 55468
rect 75740 55412 75796 55422
rect 75516 55074 75572 55086
rect 75516 55022 75518 55074
rect 75570 55022 75572 55074
rect 75404 54402 75460 54414
rect 75404 54350 75406 54402
rect 75458 54350 75460 54402
rect 75404 53956 75460 54350
rect 75404 53890 75460 53900
rect 75516 53284 75572 55022
rect 75292 53228 75572 53284
rect 75292 53172 75348 53228
rect 75292 53040 75348 53116
rect 75740 53170 75796 55356
rect 75852 54628 75908 54638
rect 75852 53842 75908 54572
rect 75852 53790 75854 53842
rect 75906 53790 75908 53842
rect 75852 53778 75908 53790
rect 75740 53118 75742 53170
rect 75794 53118 75796 53170
rect 75740 52948 75796 53118
rect 75180 52892 75460 52948
rect 75404 52612 75460 52892
rect 75292 52556 75460 52612
rect 74284 49922 74340 49934
rect 74284 49870 74286 49922
rect 74338 49870 74340 49922
rect 74284 48468 74340 49870
rect 74620 49922 74676 50540
rect 74620 49870 74622 49922
rect 74674 49870 74676 49922
rect 74620 49858 74676 49870
rect 74732 51772 74900 51828
rect 74956 52052 75012 52062
rect 74732 49700 74788 51772
rect 74956 50594 75012 51996
rect 75068 51938 75124 51950
rect 75068 51886 75070 51938
rect 75122 51886 75124 51938
rect 75068 51604 75124 51886
rect 75068 51538 75124 51548
rect 75068 51266 75124 51278
rect 75068 51214 75070 51266
rect 75122 51214 75124 51266
rect 75068 51156 75124 51214
rect 75068 51090 75124 51100
rect 74956 50542 74958 50594
rect 75010 50542 75012 50594
rect 74956 50484 75012 50542
rect 74956 50418 75012 50428
rect 75180 50372 75236 50382
rect 74284 48402 74340 48412
rect 74620 49644 74788 49700
rect 75068 50316 75180 50372
rect 74396 44436 74452 44446
rect 74396 44342 74452 44380
rect 74172 43652 74340 43708
rect 73948 41972 74004 41982
rect 73724 41970 74004 41972
rect 73724 41918 73950 41970
rect 74002 41918 74004 41970
rect 73724 41916 74004 41918
rect 73612 41804 73780 41860
rect 72716 41580 73108 41636
rect 72716 41298 72772 41580
rect 72716 41246 72718 41298
rect 72770 41246 72772 41298
rect 72716 41188 72772 41246
rect 72716 41122 72772 41132
rect 73500 40962 73556 40974
rect 73500 40910 73502 40962
rect 73554 40910 73556 40962
rect 73388 40516 73444 40526
rect 72716 40514 73444 40516
rect 72716 40462 73390 40514
rect 73442 40462 73444 40514
rect 72716 40460 73444 40462
rect 72716 39730 72772 40460
rect 73388 40450 73444 40460
rect 73500 40404 73556 40910
rect 73612 40404 73668 40414
rect 73500 40402 73668 40404
rect 73500 40350 73614 40402
rect 73666 40350 73668 40402
rect 73500 40348 73668 40350
rect 73612 40338 73668 40348
rect 72716 39678 72718 39730
rect 72770 39678 72772 39730
rect 72716 39666 72772 39678
rect 71652 36316 71876 36372
rect 72492 38612 72660 38668
rect 71596 36278 71652 36316
rect 72492 35924 72548 38612
rect 73388 36932 73444 36942
rect 73388 36594 73444 36876
rect 73388 36542 73390 36594
rect 73442 36542 73444 36594
rect 73388 36530 73444 36542
rect 73724 36036 73780 41804
rect 73836 41186 73892 41198
rect 73836 41134 73838 41186
rect 73890 41134 73892 41186
rect 73836 39732 73892 41134
rect 73948 40516 74004 41916
rect 74060 41412 74116 41422
rect 74060 41074 74116 41356
rect 74060 41022 74062 41074
rect 74114 41022 74116 41074
rect 74060 40628 74116 41022
rect 74172 40628 74228 40638
rect 74060 40626 74228 40628
rect 74060 40574 74174 40626
rect 74226 40574 74228 40626
rect 74060 40572 74228 40574
rect 74172 40562 74228 40572
rect 73948 40450 74004 40460
rect 73836 39666 73892 39676
rect 74172 37492 74228 37502
rect 74284 37492 74340 43652
rect 74620 43540 74676 49644
rect 75068 49588 75124 50316
rect 75180 50240 75236 50316
rect 75068 49522 75124 49532
rect 75180 50148 75236 50158
rect 75180 49922 75236 50092
rect 75180 49870 75182 49922
rect 75234 49870 75236 49922
rect 75180 49140 75236 49870
rect 75180 49074 75236 49084
rect 74732 47348 74788 47358
rect 74732 45330 74788 47292
rect 75068 46788 75124 46798
rect 75068 46694 75124 46732
rect 75292 46004 75348 52556
rect 75740 52162 75796 52892
rect 75740 52110 75742 52162
rect 75794 52110 75796 52162
rect 75740 52098 75796 52110
rect 75516 51940 75572 51950
rect 75516 51602 75572 51884
rect 75516 51550 75518 51602
rect 75570 51550 75572 51602
rect 75516 51538 75572 51550
rect 75852 51492 75908 51502
rect 75852 51490 76020 51492
rect 75852 51438 75854 51490
rect 75906 51438 76020 51490
rect 75852 51436 76020 51438
rect 75852 51426 75908 51436
rect 75852 50596 75908 50606
rect 75852 50502 75908 50540
rect 75964 50148 76020 51436
rect 75964 50082 76020 50092
rect 75628 50036 75684 50046
rect 75516 49924 75572 49934
rect 75516 49830 75572 49868
rect 75404 48804 75460 48814
rect 75404 48710 75460 48748
rect 74732 45278 74734 45330
rect 74786 45278 74788 45330
rect 74732 45266 74788 45278
rect 75068 46002 75348 46004
rect 75068 45950 75294 46002
rect 75346 45950 75348 46002
rect 75068 45948 75348 45950
rect 75068 45330 75124 45948
rect 75292 45938 75348 45948
rect 75404 48580 75460 48590
rect 75068 45278 75070 45330
rect 75122 45278 75124 45330
rect 75068 44660 75124 45278
rect 75068 44594 75124 44604
rect 75292 43650 75348 43662
rect 75292 43598 75294 43650
rect 75346 43598 75348 43650
rect 75180 43540 75236 43550
rect 74620 43538 75236 43540
rect 74620 43486 74622 43538
rect 74674 43486 75182 43538
rect 75234 43486 75236 43538
rect 74620 43484 75236 43486
rect 74620 43474 74676 43484
rect 75180 43474 75236 43484
rect 75180 42532 75236 42542
rect 75180 42438 75236 42476
rect 74732 41858 74788 41870
rect 74732 41806 74734 41858
rect 74786 41806 74788 41858
rect 74620 41188 74676 41198
rect 74620 41074 74676 41132
rect 74620 41022 74622 41074
rect 74674 41022 74676 41074
rect 74620 40626 74676 41022
rect 74732 41076 74788 41806
rect 75292 41748 75348 43598
rect 75292 41188 75348 41692
rect 75292 41122 75348 41132
rect 74732 41010 74788 41020
rect 75292 40964 75348 40974
rect 75292 40870 75348 40908
rect 74620 40574 74622 40626
rect 74674 40574 74676 40626
rect 74620 40562 74676 40574
rect 74844 39732 74900 39742
rect 74844 39638 74900 39676
rect 75180 39732 75236 39742
rect 74844 38948 74900 38958
rect 74844 38854 74900 38892
rect 74620 38836 74676 38846
rect 74956 38836 75012 38846
rect 74620 38834 74788 38836
rect 74620 38782 74622 38834
rect 74674 38782 74788 38834
rect 74620 38780 74788 38782
rect 74620 38770 74676 38780
rect 74732 37604 74788 38780
rect 74844 38276 74900 38286
rect 74956 38276 75012 38780
rect 74844 38274 75012 38276
rect 74844 38222 74846 38274
rect 74898 38222 75012 38274
rect 74844 38220 75012 38222
rect 75180 38274 75236 39676
rect 75180 38222 75182 38274
rect 75234 38222 75236 38274
rect 74844 38210 74900 38220
rect 75180 38210 75236 38222
rect 75404 39620 75460 48524
rect 75628 47684 75684 49980
rect 76076 49924 76132 56924
rect 76188 56978 76468 56980
rect 76188 56926 76414 56978
rect 76466 56926 76468 56978
rect 76188 56924 76468 56926
rect 76188 56084 76244 56924
rect 76412 56914 76468 56924
rect 76300 56532 76356 56542
rect 76300 56194 76356 56476
rect 76300 56142 76302 56194
rect 76354 56142 76356 56194
rect 76300 56130 76356 56142
rect 76188 54628 76244 56028
rect 76412 56084 76468 56094
rect 76412 54852 76468 56028
rect 76524 55412 76580 57596
rect 77196 56642 77252 58156
rect 77308 57092 77364 58270
rect 77532 58324 77588 59612
rect 78092 59330 78148 59948
rect 78316 62132 78596 62188
rect 78876 62242 78932 62254
rect 78876 62190 78878 62242
rect 78930 62190 78932 62242
rect 78204 59890 78260 59902
rect 78204 59838 78206 59890
rect 78258 59838 78260 59890
rect 78204 59780 78260 59838
rect 78204 59714 78260 59724
rect 78092 59278 78094 59330
rect 78146 59278 78148 59330
rect 78092 59266 78148 59278
rect 78204 59106 78260 59118
rect 78204 59054 78206 59106
rect 78258 59054 78260 59106
rect 78204 58548 78260 59054
rect 78316 58996 78372 62132
rect 78876 62020 78932 62190
rect 78876 61954 78932 61964
rect 78988 61796 79044 63870
rect 79212 63252 79268 64316
rect 79324 64306 79380 64316
rect 79324 64148 79380 64158
rect 79324 64054 79380 64092
rect 79212 63186 79268 63196
rect 79324 63364 79380 63374
rect 79324 63250 79380 63308
rect 79324 63198 79326 63250
rect 79378 63198 79380 63250
rect 78540 61740 79044 61796
rect 79100 62468 79156 62478
rect 78540 61570 78596 61740
rect 78540 61518 78542 61570
rect 78594 61518 78596 61570
rect 78428 59892 78484 59902
rect 78540 59892 78596 61518
rect 78988 61570 79044 61582
rect 78988 61518 78990 61570
rect 79042 61518 79044 61570
rect 78988 61460 79044 61518
rect 78988 61394 79044 61404
rect 78876 61012 78932 61022
rect 78764 60788 78820 60798
rect 78764 60694 78820 60732
rect 78484 59890 78596 59892
rect 78484 59838 78542 59890
rect 78594 59838 78596 59890
rect 78484 59836 78596 59838
rect 78428 59218 78484 59836
rect 78540 59826 78596 59836
rect 78428 59166 78430 59218
rect 78482 59166 78484 59218
rect 78428 59154 78484 59166
rect 78316 58940 78484 58996
rect 78204 58482 78260 58492
rect 78316 58772 78372 58782
rect 77644 58324 77700 58334
rect 77532 58268 77644 58324
rect 77644 58192 77700 58268
rect 78204 58324 78260 58334
rect 78204 58230 78260 58268
rect 78316 58322 78372 58716
rect 78316 58270 78318 58322
rect 78370 58270 78372 58322
rect 77420 58100 77476 58110
rect 77420 57874 77476 58044
rect 77420 57822 77422 57874
rect 77474 57822 77476 57874
rect 77420 57810 77476 57822
rect 77868 57540 77924 57550
rect 77756 57538 77924 57540
rect 77756 57486 77870 57538
rect 77922 57486 77924 57538
rect 77756 57484 77924 57486
rect 77308 57026 77364 57036
rect 77420 57204 77476 57214
rect 77420 56868 77476 57148
rect 77196 56590 77198 56642
rect 77250 56590 77252 56642
rect 77196 56420 77252 56590
rect 76524 55346 76580 55356
rect 76636 56194 76692 56206
rect 76636 56142 76638 56194
rect 76690 56142 76692 56194
rect 76524 55188 76580 55198
rect 76524 55094 76580 55132
rect 76188 54562 76244 54572
rect 76300 54796 76468 54852
rect 76300 53730 76356 54796
rect 76412 54628 76468 54638
rect 76412 54534 76468 54572
rect 76636 53844 76692 56142
rect 77084 56084 77140 56094
rect 77084 55990 77140 56028
rect 77196 55860 77252 56364
rect 76972 55804 77252 55860
rect 77308 56812 77476 56868
rect 77308 56306 77364 56812
rect 77308 56254 77310 56306
rect 77362 56254 77364 56306
rect 76748 54628 76804 54638
rect 76748 54534 76804 54572
rect 76636 53788 76804 53844
rect 76300 53678 76302 53730
rect 76354 53678 76356 53730
rect 76300 53666 76356 53678
rect 76412 53732 76468 53742
rect 76412 53618 76468 53676
rect 76412 53566 76414 53618
rect 76466 53566 76468 53618
rect 76412 53554 76468 53566
rect 76636 53620 76692 53630
rect 76636 53526 76692 53564
rect 76748 52948 76804 53788
rect 76748 52882 76804 52892
rect 76860 52276 76916 52286
rect 76300 52162 76356 52174
rect 76300 52110 76302 52162
rect 76354 52110 76356 52162
rect 76300 50428 76356 52110
rect 76860 51602 76916 52220
rect 76860 51550 76862 51602
rect 76914 51550 76916 51602
rect 76860 51538 76916 51550
rect 76748 51378 76804 51390
rect 76748 51326 76750 51378
rect 76802 51326 76804 51378
rect 76188 50370 76244 50382
rect 76300 50372 76580 50428
rect 76188 50318 76190 50370
rect 76242 50318 76244 50370
rect 76188 50260 76244 50318
rect 76188 50194 76244 50204
rect 76412 50036 76468 50046
rect 76412 49942 76468 49980
rect 75740 49922 76356 49924
rect 75740 49870 76078 49922
rect 76130 49870 76356 49922
rect 75740 49868 76356 49870
rect 75740 49026 75796 49868
rect 76076 49858 76132 49868
rect 76188 49140 76244 49150
rect 76188 49046 76244 49084
rect 75740 48974 75742 49026
rect 75794 48974 75796 49026
rect 75740 48962 75796 48974
rect 75516 47628 75684 47684
rect 75964 48130 76020 48142
rect 75964 48078 75966 48130
rect 76018 48078 76020 48130
rect 75516 46788 75572 47628
rect 75852 47572 75908 47582
rect 75628 47570 75908 47572
rect 75628 47518 75854 47570
rect 75906 47518 75908 47570
rect 75628 47516 75908 47518
rect 75628 46898 75684 47516
rect 75852 47506 75908 47516
rect 75628 46846 75630 46898
rect 75682 46846 75684 46898
rect 75628 46834 75684 46846
rect 75852 46900 75908 46910
rect 75852 46806 75908 46844
rect 75516 46656 75572 46732
rect 75964 46452 76020 48078
rect 76300 47572 76356 49868
rect 76524 48692 76580 50372
rect 76748 50372 76804 51326
rect 76748 50306 76804 50316
rect 76860 50484 76916 50494
rect 76860 50034 76916 50428
rect 76860 49982 76862 50034
rect 76914 49982 76916 50034
rect 76860 49970 76916 49982
rect 76972 49252 77028 55804
rect 77196 55188 77252 55198
rect 77196 55094 77252 55132
rect 77308 53172 77364 56254
rect 77420 56644 77476 56654
rect 77420 56194 77476 56588
rect 77420 56142 77422 56194
rect 77474 56142 77476 56194
rect 77420 56130 77476 56142
rect 77644 56642 77700 56654
rect 77644 56590 77646 56642
rect 77698 56590 77700 56642
rect 77644 55300 77700 56590
rect 77756 56308 77812 57484
rect 77868 57474 77924 57484
rect 78316 57204 78372 58270
rect 78428 58548 78484 58940
rect 78428 57876 78484 58492
rect 78876 58546 78932 60956
rect 78988 59332 79044 59342
rect 78988 59238 79044 59276
rect 78876 58494 78878 58546
rect 78930 58494 78932 58546
rect 78540 58212 78596 58222
rect 78540 58118 78596 58156
rect 78876 58100 78932 58494
rect 79100 58436 79156 62412
rect 79324 61124 79380 63198
rect 79436 62468 79492 64988
rect 79660 64148 79716 65100
rect 79660 64082 79716 64092
rect 79660 63700 79716 63710
rect 79660 63140 79716 63644
rect 79548 63138 79716 63140
rect 79548 63086 79662 63138
rect 79714 63086 79716 63138
rect 79548 63084 79716 63086
rect 79548 62916 79604 63084
rect 79660 63074 79716 63084
rect 79772 62916 79828 65436
rect 79996 65398 80052 65436
rect 80108 65380 80164 65390
rect 79996 64708 80052 64718
rect 79996 64614 80052 64652
rect 79884 64260 79940 64270
rect 79884 64146 79940 64204
rect 79884 64094 79886 64146
rect 79938 64094 79940 64146
rect 79884 64082 79940 64094
rect 79996 64036 80052 64046
rect 79548 62850 79604 62860
rect 79660 62860 79828 62916
rect 79884 63812 79940 63822
rect 79436 62336 79492 62412
rect 79660 62020 79716 62860
rect 79772 62466 79828 62478
rect 79772 62414 79774 62466
rect 79826 62414 79828 62466
rect 79772 62244 79828 62414
rect 79772 62178 79828 62188
rect 79660 61954 79716 61964
rect 79884 61796 79940 63756
rect 79772 61740 79940 61796
rect 79548 61460 79604 61470
rect 79212 61068 79380 61124
rect 79436 61458 79604 61460
rect 79436 61406 79550 61458
rect 79602 61406 79604 61458
rect 79436 61404 79604 61406
rect 79436 61348 79492 61404
rect 79548 61394 79604 61404
rect 79212 60564 79268 61068
rect 79324 60900 79380 60910
rect 79324 60806 79380 60844
rect 79436 60676 79492 61292
rect 79660 61348 79716 61358
rect 79660 61254 79716 61292
rect 79660 61012 79716 61022
rect 79660 60898 79716 60956
rect 79660 60846 79662 60898
rect 79714 60846 79716 60898
rect 79660 60834 79716 60846
rect 79436 60620 79716 60676
rect 79212 60508 79604 60564
rect 79436 59892 79492 59902
rect 79100 58370 79156 58380
rect 79212 59890 79492 59892
rect 79212 59838 79438 59890
rect 79490 59838 79492 59890
rect 79212 59836 79492 59838
rect 78876 58034 78932 58044
rect 78428 57810 78484 57820
rect 78540 57988 78596 57998
rect 78540 57762 78596 57932
rect 78876 57876 78932 57886
rect 78876 57782 78932 57820
rect 78540 57710 78542 57762
rect 78594 57710 78596 57762
rect 78540 57698 78596 57710
rect 78316 57138 78372 57148
rect 78988 56980 79044 56990
rect 78988 56886 79044 56924
rect 78204 56866 78260 56878
rect 78204 56814 78206 56866
rect 78258 56814 78260 56866
rect 77756 56242 77812 56252
rect 77868 56532 77924 56542
rect 77868 56306 77924 56476
rect 77868 56254 77870 56306
rect 77922 56254 77924 56306
rect 77868 56242 77924 56254
rect 77756 55300 77812 55310
rect 77644 55298 77812 55300
rect 77644 55246 77758 55298
rect 77810 55246 77812 55298
rect 77644 55244 77812 55246
rect 77644 54740 77700 55244
rect 77756 55234 77812 55244
rect 78204 55300 78260 56814
rect 78876 56194 78932 56206
rect 78876 56142 78878 56194
rect 78930 56142 78932 56194
rect 78764 56082 78820 56094
rect 78764 56030 78766 56082
rect 78818 56030 78820 56082
rect 78428 55860 78484 55870
rect 78204 55234 78260 55244
rect 78316 55298 78372 55310
rect 78316 55246 78318 55298
rect 78370 55246 78372 55298
rect 77644 54674 77700 54684
rect 77756 54516 77812 54526
rect 77532 54460 77756 54516
rect 77420 53732 77476 53742
rect 77532 53732 77588 54460
rect 77756 54422 77812 54460
rect 77420 53730 77588 53732
rect 77420 53678 77422 53730
rect 77474 53678 77588 53730
rect 77420 53676 77588 53678
rect 77420 53666 77476 53676
rect 77308 53106 77364 53116
rect 77196 51938 77252 51950
rect 77196 51886 77198 51938
rect 77250 51886 77252 51938
rect 77084 51380 77140 51390
rect 77084 51286 77140 51324
rect 77196 51156 77252 51886
rect 77420 51940 77476 51950
rect 77420 51602 77476 51884
rect 77420 51550 77422 51602
rect 77474 51550 77476 51602
rect 77420 51538 77476 51550
rect 77084 51100 77252 51156
rect 77084 50372 77140 51100
rect 77084 50306 77140 50316
rect 77196 50484 77252 50560
rect 76524 48626 76580 48636
rect 76860 49196 77028 49252
rect 76524 48468 76580 48478
rect 76412 47572 76468 47582
rect 76300 47570 76468 47572
rect 76300 47518 76414 47570
rect 76466 47518 76468 47570
rect 76300 47516 76468 47518
rect 76412 47460 76468 47516
rect 76412 47394 76468 47404
rect 76300 46900 76356 46910
rect 76300 46786 76356 46844
rect 76412 46900 76468 46910
rect 76524 46900 76580 48412
rect 76748 48244 76804 48254
rect 76748 48150 76804 48188
rect 76412 46898 76580 46900
rect 76412 46846 76414 46898
rect 76466 46846 76580 46898
rect 76412 46844 76580 46846
rect 76412 46834 76468 46844
rect 76300 46734 76302 46786
rect 76354 46734 76356 46786
rect 76300 46722 76356 46734
rect 76412 46452 76468 46462
rect 75964 46450 76468 46452
rect 75964 46398 76414 46450
rect 76466 46398 76468 46450
rect 75964 46396 76468 46398
rect 76412 46386 76468 46396
rect 76076 46004 76132 46014
rect 76076 45910 76132 45948
rect 75628 45218 75684 45230
rect 75628 45166 75630 45218
rect 75682 45166 75684 45218
rect 75628 44436 75684 45166
rect 75964 45108 76020 45118
rect 75964 45106 76356 45108
rect 75964 45054 75966 45106
rect 76018 45054 76356 45106
rect 75964 45052 76356 45054
rect 75964 45042 76020 45052
rect 76076 44660 76132 44670
rect 75628 44370 75684 44380
rect 75964 44436 76020 44446
rect 75964 43538 76020 44380
rect 75964 43486 75966 43538
rect 76018 43486 76020 43538
rect 75964 43474 76020 43486
rect 75740 42756 75796 42766
rect 75740 42662 75796 42700
rect 75852 41300 75908 41310
rect 75852 41206 75908 41244
rect 74732 37548 75348 37604
rect 73948 37490 74340 37492
rect 73948 37438 74174 37490
rect 74226 37438 74340 37490
rect 73948 37436 74340 37438
rect 75292 37490 75348 37548
rect 75292 37438 75294 37490
rect 75346 37438 75348 37490
rect 73388 35980 73780 36036
rect 73836 36484 73892 36494
rect 73948 36484 74004 37436
rect 74172 37426 74228 37436
rect 75292 37426 75348 37438
rect 74620 37154 74676 37166
rect 74620 37102 74622 37154
rect 74674 37102 74676 37154
rect 73836 36482 74004 36484
rect 73836 36430 73838 36482
rect 73890 36430 74004 36482
rect 73836 36428 74004 36430
rect 74060 36932 74116 36942
rect 72492 35868 72772 35924
rect 71708 35810 71764 35822
rect 71708 35758 71710 35810
rect 71762 35758 71764 35810
rect 71148 34802 71204 34814
rect 71148 34750 71150 34802
rect 71202 34750 71204 34802
rect 70812 34692 70868 34702
rect 70476 34690 70868 34692
rect 70476 34638 70814 34690
rect 70866 34638 70868 34690
rect 70476 34636 70868 34638
rect 70476 33458 70532 34636
rect 70812 34626 70868 34636
rect 71148 34356 71204 34750
rect 71148 34290 71204 34300
rect 70476 33406 70478 33458
rect 70530 33406 70532 33458
rect 70476 33394 70532 33406
rect 70812 33348 70868 33358
rect 70252 32674 70308 33068
rect 70252 32622 70254 32674
rect 70306 32622 70308 32674
rect 69580 32452 69636 32462
rect 69580 32358 69636 32396
rect 69244 32340 69300 32350
rect 69244 32246 69300 32284
rect 70252 31892 70308 32622
rect 70364 33236 70420 33246
rect 70364 32562 70420 33180
rect 70364 32510 70366 32562
rect 70418 32510 70420 32562
rect 70364 32498 70420 32510
rect 70812 32564 70868 33292
rect 71372 33236 71428 33246
rect 71372 32786 71428 33180
rect 71372 32734 71374 32786
rect 71426 32734 71428 32786
rect 71372 32722 71428 32734
rect 70924 32564 70980 32574
rect 70812 32508 70924 32564
rect 70364 31892 70420 31902
rect 68572 31890 68740 31892
rect 68572 31838 68574 31890
rect 68626 31838 68740 31890
rect 68572 31836 68740 31838
rect 69692 31890 70420 31892
rect 69692 31838 70366 31890
rect 70418 31838 70420 31890
rect 69692 31836 70420 31838
rect 68572 31826 68628 31836
rect 68012 31726 68014 31778
rect 68066 31726 68068 31778
rect 68012 31714 68068 31726
rect 69356 31780 69412 31790
rect 66668 31614 66670 31666
rect 66722 31614 66724 31666
rect 66668 31602 66724 31614
rect 67676 31668 67732 31678
rect 67676 31574 67732 31612
rect 69356 31666 69412 31724
rect 69356 31614 69358 31666
rect 69410 31614 69412 31666
rect 57372 31502 57374 31554
rect 57426 31502 57428 31554
rect 56028 3444 56084 3454
rect 56140 3444 56196 3454
rect 56028 3442 56140 3444
rect 56028 3390 56030 3442
rect 56082 3390 56140 3442
rect 56028 3388 56140 3390
rect 56028 3378 56084 3388
rect 54348 3266 54404 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 45276 2706 45332 2716
rect 56140 800 56196 3388
rect 56700 3444 56756 3454
rect 56700 3350 56756 3388
rect 57036 3330 57092 3342
rect 57036 3278 57038 3330
rect 57090 3278 57092 3330
rect 57036 2996 57092 3278
rect 57036 2930 57092 2940
rect 57372 2884 57428 31502
rect 69020 30884 69076 30894
rect 69356 30884 69412 31614
rect 69692 31666 69748 31836
rect 70364 31826 70420 31836
rect 69692 31614 69694 31666
rect 69746 31614 69748 31666
rect 69692 31602 69748 31614
rect 70812 31778 70868 32508
rect 70924 32432 70980 32508
rect 71708 31948 71764 35758
rect 71932 35698 71988 35710
rect 71932 35646 71934 35698
rect 71986 35646 71988 35698
rect 71820 35140 71876 35150
rect 71932 35140 71988 35646
rect 72604 35588 72660 35598
rect 71820 35138 71988 35140
rect 71820 35086 71822 35138
rect 71874 35086 71988 35138
rect 71820 35084 71988 35086
rect 72380 35586 72660 35588
rect 72380 35534 72606 35586
rect 72658 35534 72660 35586
rect 72380 35532 72660 35534
rect 71820 35074 71876 35084
rect 72380 35028 72436 35532
rect 72604 35522 72660 35532
rect 72156 34916 72212 34926
rect 72156 34822 72212 34860
rect 72380 34802 72436 34972
rect 72380 34750 72382 34802
rect 72434 34750 72436 34802
rect 72380 34738 72436 34750
rect 72604 34916 72660 34926
rect 72044 34692 72100 34702
rect 72044 32562 72100 34636
rect 72604 34132 72660 34860
rect 72716 34804 72772 35868
rect 72716 34802 72884 34804
rect 72716 34750 72718 34802
rect 72770 34750 72884 34802
rect 72716 34748 72884 34750
rect 72716 34738 72772 34748
rect 72604 33458 72660 34076
rect 72828 33570 72884 34748
rect 72828 33518 72830 33570
rect 72882 33518 72884 33570
rect 72828 33506 72884 33518
rect 72604 33406 72606 33458
rect 72658 33406 72660 33458
rect 72604 33394 72660 33406
rect 73052 33124 73108 33134
rect 73052 33030 73108 33068
rect 72604 32788 72660 32798
rect 72604 32694 72660 32732
rect 72044 32510 72046 32562
rect 72098 32510 72100 32562
rect 72044 32498 72100 32510
rect 73276 32564 73332 32574
rect 73276 32470 73332 32508
rect 71596 31892 71764 31948
rect 71596 31890 71652 31892
rect 71596 31838 71598 31890
rect 71650 31838 71652 31890
rect 71596 31826 71652 31838
rect 70812 31726 70814 31778
rect 70866 31726 70868 31778
rect 70588 31220 70644 31230
rect 70812 31220 70868 31726
rect 70588 31218 70868 31220
rect 70588 31166 70590 31218
rect 70642 31166 70868 31218
rect 70588 31164 70868 31166
rect 70588 31154 70644 31164
rect 69020 30882 69412 30884
rect 69020 30830 69022 30882
rect 69074 30830 69412 30882
rect 69020 30828 69412 30830
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 67788 3444 67844 3454
rect 67788 3350 67844 3388
rect 68796 3444 68852 3454
rect 57372 2818 57428 2828
rect 68796 2324 68852 3388
rect 69020 2772 69076 30828
rect 73388 12740 73444 35980
rect 73500 35586 73556 35598
rect 73500 35534 73502 35586
rect 73554 35534 73556 35586
rect 73500 35028 73556 35534
rect 73500 34962 73556 34972
rect 73724 34916 73780 34926
rect 73724 34822 73780 34860
rect 73500 34356 73556 34366
rect 73836 34356 73892 36428
rect 74060 35922 74116 36876
rect 74620 36932 74676 37102
rect 74620 36866 74676 36876
rect 75404 36932 75460 39564
rect 75516 40516 75572 40526
rect 75516 38834 75572 40460
rect 75852 39732 75908 39742
rect 75516 38782 75518 38834
rect 75570 38782 75572 38834
rect 75516 38770 75572 38782
rect 75740 39730 75908 39732
rect 75740 39678 75854 39730
rect 75906 39678 75908 39730
rect 75740 39676 75908 39678
rect 75628 38724 75684 38734
rect 75628 37266 75684 38668
rect 75740 37380 75796 39676
rect 75852 39666 75908 39676
rect 75852 38052 75908 38062
rect 75852 37958 75908 37996
rect 75964 37940 76020 37950
rect 75964 37846 76020 37884
rect 75852 37380 75908 37390
rect 75740 37324 75852 37380
rect 75852 37286 75908 37324
rect 75628 37214 75630 37266
rect 75682 37214 75684 37266
rect 75628 37202 75684 37214
rect 74060 35870 74062 35922
rect 74114 35870 74116 35922
rect 74060 35858 74116 35870
rect 74284 36594 74340 36606
rect 74284 36542 74286 36594
rect 74338 36542 74340 36594
rect 74284 35924 74340 36542
rect 74284 35858 74340 35868
rect 74620 36484 74676 36494
rect 74396 35812 74452 35822
rect 74396 35026 74452 35756
rect 74396 34974 74398 35026
rect 74450 34974 74452 35026
rect 74396 34962 74452 34974
rect 73500 34262 73556 34300
rect 73724 34300 73892 34356
rect 73500 33570 73556 33582
rect 73500 33518 73502 33570
rect 73554 33518 73556 33570
rect 73500 33458 73556 33518
rect 73500 33406 73502 33458
rect 73554 33406 73556 33458
rect 73500 31948 73556 33406
rect 73724 33348 73780 34300
rect 74396 34242 74452 34254
rect 74396 34190 74398 34242
rect 74450 34190 74452 34242
rect 73836 34132 73892 34142
rect 73836 34038 73892 34076
rect 74396 33908 74452 34190
rect 74620 34132 74676 36428
rect 74956 36484 75012 36494
rect 74956 36390 75012 36428
rect 75404 36482 75460 36876
rect 75404 36430 75406 36482
rect 75458 36430 75460 36482
rect 75404 36418 75460 36430
rect 76076 36596 76132 44604
rect 76300 43762 76356 45052
rect 76748 45106 76804 45118
rect 76748 45054 76750 45106
rect 76802 45054 76804 45106
rect 76524 44436 76580 44446
rect 76524 44342 76580 44380
rect 76300 43710 76302 43762
rect 76354 43710 76356 43762
rect 76300 43698 76356 43710
rect 76748 42980 76804 45054
rect 76748 42914 76804 42924
rect 76188 42532 76244 42542
rect 76188 42438 76244 42476
rect 76860 42420 76916 49196
rect 77196 49028 77252 50428
rect 77532 49810 77588 53676
rect 78092 53620 78148 53630
rect 78092 53526 78148 53564
rect 77644 53172 77700 53182
rect 78316 53172 78372 55246
rect 78428 54626 78484 55804
rect 78428 54574 78430 54626
rect 78482 54574 78484 54626
rect 78428 54562 78484 54574
rect 78764 53732 78820 56030
rect 78876 56084 78932 56142
rect 78876 56028 79044 56084
rect 78876 55860 78932 55870
rect 78876 55766 78932 55804
rect 78988 55522 79044 56028
rect 78988 55470 78990 55522
rect 79042 55470 79044 55522
rect 78988 55458 79044 55470
rect 79212 55412 79268 59836
rect 79436 59826 79492 59836
rect 79324 59220 79380 59230
rect 79324 59126 79380 59164
rect 79324 58210 79380 58222
rect 79324 58158 79326 58210
rect 79378 58158 79380 58210
rect 79324 58100 79380 58158
rect 79324 57764 79380 58044
rect 79324 57698 79380 57708
rect 79436 58212 79492 58222
rect 79436 57762 79492 58156
rect 79548 57988 79604 60508
rect 79660 58212 79716 60620
rect 79772 60116 79828 61740
rect 79884 61572 79940 61582
rect 79996 61572 80052 63980
rect 80108 63138 80164 65324
rect 80332 65378 80388 65390
rect 80332 65326 80334 65378
rect 80386 65326 80388 65378
rect 80332 65044 80388 65326
rect 80332 64978 80388 64988
rect 80220 64484 80276 64494
rect 80220 64482 80612 64484
rect 80220 64430 80222 64482
rect 80274 64430 80612 64482
rect 80220 64428 80612 64430
rect 80220 64418 80276 64428
rect 80220 64148 80276 64158
rect 80220 64034 80276 64092
rect 80220 63982 80222 64034
rect 80274 63982 80276 64034
rect 80220 63970 80276 63982
rect 80108 63086 80110 63138
rect 80162 63086 80164 63138
rect 80108 63074 80164 63086
rect 80444 63924 80500 63934
rect 80332 62914 80388 62926
rect 80332 62862 80334 62914
rect 80386 62862 80388 62914
rect 80332 62468 80388 62862
rect 80332 62402 80388 62412
rect 80220 62242 80276 62254
rect 80220 62190 80222 62242
rect 80274 62190 80276 62242
rect 79884 61570 80052 61572
rect 79884 61518 79886 61570
rect 79938 61518 80052 61570
rect 79884 61516 80052 61518
rect 80108 62020 80164 62030
rect 79884 61506 79940 61516
rect 79772 60002 79828 60060
rect 79772 59950 79774 60002
rect 79826 59950 79828 60002
rect 79772 59938 79828 59950
rect 79996 60452 80052 60462
rect 79996 59668 80052 60396
rect 80108 60004 80164 61964
rect 80220 61908 80276 62190
rect 80220 61842 80276 61852
rect 80444 61682 80500 63868
rect 80556 62580 80612 64428
rect 80668 64372 80724 65884
rect 80780 66388 80836 66398
rect 80780 64706 80836 66332
rect 81452 66386 81508 67118
rect 81564 67060 81620 67070
rect 81564 66966 81620 67004
rect 81452 66334 81454 66386
rect 81506 66334 81508 66386
rect 81452 66052 81508 66334
rect 81116 65996 81508 66052
rect 81004 65828 81060 65838
rect 80780 64654 80782 64706
rect 80834 64654 80836 64706
rect 80780 64642 80836 64654
rect 80892 65716 80948 65726
rect 80892 64594 80948 65660
rect 81004 65604 81060 65772
rect 81004 65538 81060 65548
rect 81116 65380 81172 65996
rect 81276 65884 81540 65894
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81276 65818 81540 65828
rect 81116 65314 81172 65324
rect 81228 65378 81284 65390
rect 81228 65326 81230 65378
rect 81282 65326 81284 65378
rect 81228 65044 81284 65326
rect 81228 64978 81284 64988
rect 81564 64930 81620 64942
rect 81564 64878 81566 64930
rect 81618 64878 81620 64930
rect 81564 64818 81620 64878
rect 81564 64766 81566 64818
rect 81618 64766 81620 64818
rect 81564 64754 81620 64766
rect 80892 64542 80894 64594
rect 80946 64542 80948 64594
rect 80892 64530 80948 64542
rect 81004 64596 81060 64606
rect 80668 64316 80948 64372
rect 80556 62514 80612 62524
rect 80668 63252 80724 63262
rect 80668 62916 80724 63196
rect 80444 61630 80446 61682
rect 80498 61630 80500 61682
rect 80444 61618 80500 61630
rect 80668 61570 80724 62860
rect 80668 61518 80670 61570
rect 80722 61518 80724 61570
rect 80668 61506 80724 61518
rect 80780 62244 80836 62254
rect 80780 61570 80836 62188
rect 80892 62188 80948 64316
rect 81004 63138 81060 64540
rect 81116 64482 81172 64494
rect 81116 64430 81118 64482
rect 81170 64430 81172 64482
rect 81116 64148 81172 64430
rect 81276 64316 81540 64326
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81276 64250 81540 64260
rect 81116 64082 81172 64092
rect 81564 63924 81620 63934
rect 81564 63830 81620 63868
rect 81004 63086 81006 63138
rect 81058 63086 81060 63138
rect 81004 63028 81060 63086
rect 81564 63252 81620 63262
rect 81676 63252 81732 70812
rect 82796 70866 82964 70868
rect 82796 70814 82910 70866
rect 82962 70814 82964 70866
rect 82796 70812 82964 70814
rect 81900 70196 81956 70206
rect 81900 69524 81956 70140
rect 81900 69410 81956 69468
rect 81900 69358 81902 69410
rect 81954 69358 81956 69410
rect 81900 69346 81956 69358
rect 82572 70194 82628 70206
rect 82572 70142 82574 70194
rect 82626 70142 82628 70194
rect 82124 69300 82180 69310
rect 82124 69206 82180 69244
rect 82572 68964 82628 70142
rect 82684 69524 82740 69534
rect 82796 69524 82852 70812
rect 82908 70532 82964 70812
rect 82908 70466 82964 70476
rect 83020 70756 83076 70926
rect 82684 69522 82852 69524
rect 82684 69470 82686 69522
rect 82738 69470 82852 69522
rect 82684 69468 82852 69470
rect 82684 69300 82740 69468
rect 82684 69234 82740 69244
rect 83020 69076 83076 70700
rect 83244 70306 83300 73390
rect 83244 70254 83246 70306
rect 83298 70254 83300 70306
rect 83244 70242 83300 70254
rect 83356 70532 83412 70542
rect 83244 69300 83300 69310
rect 82572 68898 82628 68908
rect 82908 69020 83076 69076
rect 83132 69298 83300 69300
rect 83132 69246 83246 69298
rect 83298 69246 83300 69298
rect 83132 69244 83300 69246
rect 82572 67844 82628 67854
rect 82572 67750 82628 67788
rect 82572 67172 82628 67182
rect 82012 66946 82068 66958
rect 82012 66894 82014 66946
rect 82066 66894 82068 66946
rect 82012 66836 82068 66894
rect 82012 66770 82068 66780
rect 81900 66500 81956 66510
rect 81900 66386 81956 66444
rect 81900 66334 81902 66386
rect 81954 66334 81956 66386
rect 81900 66322 81956 66334
rect 82124 66500 82180 66510
rect 81900 65604 81956 65614
rect 81788 65378 81844 65390
rect 81788 65326 81790 65378
rect 81842 65326 81844 65378
rect 81788 64596 81844 65326
rect 81900 64818 81956 65548
rect 81900 64766 81902 64818
rect 81954 64766 81956 64818
rect 81900 64754 81956 64766
rect 81788 64530 81844 64540
rect 82124 64372 82180 66444
rect 82348 66388 82404 66398
rect 82348 66294 82404 66332
rect 82236 65378 82292 65390
rect 82236 65326 82238 65378
rect 82290 65326 82292 65378
rect 82236 65156 82292 65326
rect 82236 65090 82292 65100
rect 81900 64316 82180 64372
rect 82236 64930 82292 64942
rect 82236 64878 82238 64930
rect 82290 64878 82292 64930
rect 81900 64146 81956 64316
rect 81900 64094 81902 64146
rect 81954 64094 81956 64146
rect 81900 64082 81956 64094
rect 82012 64148 82068 64186
rect 82012 64082 82068 64092
rect 81788 63924 81844 63934
rect 82124 63924 82180 63934
rect 81788 63830 81844 63868
rect 82012 63922 82180 63924
rect 82012 63870 82126 63922
rect 82178 63870 82180 63922
rect 82012 63868 82180 63870
rect 81620 63196 81732 63252
rect 81564 63138 81620 63196
rect 81564 63086 81566 63138
rect 81618 63086 81620 63138
rect 81564 63074 81620 63086
rect 81004 62962 81060 62972
rect 82012 62916 82068 63868
rect 82124 63858 82180 63868
rect 82236 62916 82292 64878
rect 82348 64482 82404 64494
rect 82348 64430 82350 64482
rect 82402 64430 82404 64482
rect 82348 63364 82404 64430
rect 82348 63298 82404 63308
rect 82460 64260 82516 64270
rect 81676 62860 82068 62916
rect 82124 62860 82292 62916
rect 82348 63138 82404 63150
rect 82348 63086 82350 63138
rect 82402 63086 82404 63138
rect 81276 62748 81540 62758
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81276 62682 81540 62692
rect 81564 62580 81620 62590
rect 81676 62580 81732 62860
rect 81564 62578 81732 62580
rect 81564 62526 81566 62578
rect 81618 62526 81732 62578
rect 81564 62524 81732 62526
rect 81900 62580 81956 62590
rect 81564 62514 81620 62524
rect 81340 62468 81396 62478
rect 81340 62374 81396 62412
rect 81900 62466 81956 62524
rect 81900 62414 81902 62466
rect 81954 62414 81956 62466
rect 81900 62402 81956 62414
rect 81676 62356 81732 62366
rect 81676 62262 81732 62300
rect 82124 62356 82180 62860
rect 82124 62188 82180 62300
rect 80892 62132 81060 62188
rect 80780 61518 80782 61570
rect 80834 61518 80836 61570
rect 80780 61506 80836 61518
rect 80332 61458 80388 61470
rect 80332 61406 80334 61458
rect 80386 61406 80388 61458
rect 80220 60786 80276 60798
rect 80220 60734 80222 60786
rect 80274 60734 80276 60786
rect 80220 60564 80276 60734
rect 80220 60498 80276 60508
rect 80220 60004 80276 60014
rect 80108 60002 80276 60004
rect 80108 59950 80222 60002
rect 80274 59950 80276 60002
rect 80108 59948 80276 59950
rect 80220 59892 80276 59948
rect 80332 59892 80388 61406
rect 80556 60898 80612 60910
rect 80556 60846 80558 60898
rect 80610 60846 80612 60898
rect 80556 60116 80612 60846
rect 80556 60060 80948 60116
rect 80892 60002 80948 60060
rect 80892 59950 80894 60002
rect 80946 59950 80948 60002
rect 80444 59892 80500 59902
rect 80332 59890 80500 59892
rect 80332 59838 80446 59890
rect 80498 59838 80500 59890
rect 80332 59836 80500 59838
rect 80220 59826 80276 59836
rect 80444 59826 80500 59836
rect 79996 59612 80388 59668
rect 80332 59442 80388 59612
rect 80332 59390 80334 59442
rect 80386 59390 80388 59442
rect 80332 59378 80388 59390
rect 80892 59444 80948 59950
rect 80892 59378 80948 59388
rect 79996 59220 80052 59230
rect 79772 59108 79828 59118
rect 79772 59014 79828 59052
rect 79772 58436 79828 58446
rect 79772 58342 79828 58380
rect 79660 58156 79828 58212
rect 79548 57932 79716 57988
rect 79436 57710 79438 57762
rect 79490 57710 79492 57762
rect 79436 57698 79492 57710
rect 79548 57764 79604 57774
rect 79548 57670 79604 57708
rect 79548 57426 79604 57438
rect 79548 57374 79550 57426
rect 79602 57374 79604 57426
rect 79548 56980 79604 57374
rect 79548 56914 79604 56924
rect 79436 56644 79492 56654
rect 79436 56306 79492 56588
rect 79436 56254 79438 56306
rect 79490 56254 79492 56306
rect 79436 56242 79492 56254
rect 79100 55356 79268 55412
rect 79100 55300 79156 55356
rect 78988 55244 79156 55300
rect 78988 55186 79044 55244
rect 78988 55134 78990 55186
rect 79042 55134 79044 55186
rect 78988 55122 79044 55134
rect 79100 55130 79156 55142
rect 79100 55078 79102 55130
rect 79154 55078 79156 55130
rect 79100 54628 79156 55078
rect 79100 54562 79156 54572
rect 79212 54404 79268 55356
rect 79212 54338 79268 54348
rect 79548 54628 79604 54638
rect 77644 52276 77700 53116
rect 77644 52144 77700 52220
rect 77868 53116 78372 53172
rect 78428 53172 78484 53182
rect 77532 49758 77534 49810
rect 77586 49758 77588 49810
rect 77308 49028 77364 49038
rect 77196 48972 77308 49028
rect 77308 48896 77364 48972
rect 77532 48244 77588 49758
rect 77644 50372 77700 50382
rect 77644 48914 77700 50316
rect 77644 48862 77646 48914
rect 77698 48862 77700 48914
rect 77644 48850 77700 48862
rect 77756 49028 77812 49038
rect 77532 48178 77588 48188
rect 77644 48692 77700 48702
rect 77644 48242 77700 48636
rect 77644 48190 77646 48242
rect 77698 48190 77700 48242
rect 77308 48130 77364 48142
rect 77308 48078 77310 48130
rect 77362 48078 77364 48130
rect 77308 47684 77364 48078
rect 77084 47628 77364 47684
rect 76636 42364 76916 42420
rect 76972 46564 77028 46574
rect 77084 46564 77140 47628
rect 77644 47572 77700 48190
rect 77196 47460 77252 47470
rect 77644 47460 77700 47516
rect 77196 47366 77252 47404
rect 77532 47404 77700 47460
rect 77532 46898 77588 47404
rect 77644 47236 77700 47246
rect 77756 47236 77812 48972
rect 77644 47234 77812 47236
rect 77644 47182 77646 47234
rect 77698 47182 77812 47234
rect 77644 47180 77812 47182
rect 77644 47170 77700 47180
rect 77532 46846 77534 46898
rect 77586 46846 77588 46898
rect 77532 46834 77588 46846
rect 76972 46562 77140 46564
rect 76972 46510 76974 46562
rect 77026 46510 77140 46562
rect 76972 46508 77140 46510
rect 76636 41636 76692 42364
rect 76972 42308 77028 46508
rect 77420 45780 77476 45790
rect 77308 45666 77364 45678
rect 77308 45614 77310 45666
rect 77362 45614 77364 45666
rect 77084 45218 77140 45230
rect 77084 45166 77086 45218
rect 77138 45166 77140 45218
rect 77084 43652 77140 45166
rect 77084 43586 77140 43596
rect 77196 45108 77252 45118
rect 77196 43538 77252 45052
rect 77196 43486 77198 43538
rect 77250 43486 77252 43538
rect 77196 43474 77252 43486
rect 76972 42252 77140 42308
rect 77084 41972 77140 42252
rect 77308 42084 77364 45614
rect 77420 44546 77476 45724
rect 77868 45668 77924 53116
rect 78428 53078 78484 53116
rect 78652 53172 78708 53182
rect 78764 53172 78820 53676
rect 78652 53170 78820 53172
rect 78652 53118 78654 53170
rect 78706 53118 78820 53170
rect 78652 53116 78820 53118
rect 79548 53170 79604 54572
rect 79548 53118 79550 53170
rect 79602 53118 79604 53170
rect 78652 53106 78708 53116
rect 79548 53106 79604 53118
rect 78316 52948 78372 52958
rect 78316 52854 78372 52892
rect 79100 52948 79156 52958
rect 79100 52854 79156 52892
rect 78764 52612 78820 52622
rect 78764 52274 78820 52556
rect 78764 52222 78766 52274
rect 78818 52222 78820 52274
rect 78764 52210 78820 52222
rect 79100 52612 79156 52622
rect 78316 51492 78372 51502
rect 78316 51398 78372 51436
rect 79100 51490 79156 52556
rect 79100 51438 79102 51490
rect 79154 51438 79156 51490
rect 78204 51380 78260 51390
rect 78204 51286 78260 51324
rect 78316 51154 78372 51166
rect 78316 51102 78318 51154
rect 78370 51102 78372 51154
rect 78316 49922 78372 51102
rect 79100 50260 79156 51438
rect 79212 51492 79268 51502
rect 79436 51492 79492 51502
rect 79212 51490 79380 51492
rect 79212 51438 79214 51490
rect 79266 51438 79380 51490
rect 79212 51436 79380 51438
rect 79212 51426 79268 51436
rect 79324 50932 79380 51436
rect 79436 51398 79492 51436
rect 79100 50194 79156 50204
rect 79212 50876 79380 50932
rect 78764 50148 78820 50158
rect 78316 49870 78318 49922
rect 78370 49870 78372 49922
rect 78316 49858 78372 49870
rect 78428 49924 78484 49934
rect 77980 49140 78036 49150
rect 77980 46898 78036 49084
rect 78428 49140 78484 49868
rect 78428 49026 78484 49084
rect 78428 48974 78430 49026
rect 78482 48974 78484 49026
rect 78428 48962 78484 48974
rect 78652 49028 78708 49038
rect 78092 48802 78148 48814
rect 78316 48804 78372 48814
rect 78092 48750 78094 48802
rect 78146 48750 78148 48802
rect 78092 48468 78148 48750
rect 78092 48402 78148 48412
rect 78204 48802 78372 48804
rect 78204 48750 78318 48802
rect 78370 48750 78372 48802
rect 78204 48748 78372 48750
rect 78092 48244 78148 48254
rect 78204 48244 78260 48748
rect 78316 48738 78372 48748
rect 78316 48468 78372 48478
rect 78316 48374 78372 48412
rect 78092 48242 78260 48244
rect 78092 48190 78094 48242
rect 78146 48190 78260 48242
rect 78092 48188 78260 48190
rect 78652 48244 78708 48972
rect 78092 48132 78148 48188
rect 78092 48066 78148 48076
rect 78652 47570 78708 48188
rect 78652 47518 78654 47570
rect 78706 47518 78708 47570
rect 78652 47506 78708 47518
rect 78764 48354 78820 50092
rect 79212 49700 79268 50876
rect 79548 50596 79604 50606
rect 79548 50502 79604 50540
rect 79660 50428 79716 57932
rect 79772 55972 79828 58156
rect 79996 57092 80052 59164
rect 81004 58772 81060 62132
rect 81676 62132 81732 62142
rect 81452 61796 81508 61806
rect 81452 61458 81508 61740
rect 81452 61406 81454 61458
rect 81506 61406 81508 61458
rect 81452 61394 81508 61406
rect 81676 61570 81732 62076
rect 81676 61518 81678 61570
rect 81730 61518 81732 61570
rect 81276 61180 81540 61190
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81276 61114 81540 61124
rect 81676 60900 81732 61518
rect 81676 60834 81732 60844
rect 81788 62132 82180 62188
rect 82236 62692 82292 62702
rect 81340 60786 81396 60798
rect 81340 60734 81342 60786
rect 81394 60734 81396 60786
rect 81340 60228 81396 60734
rect 81452 60564 81508 60574
rect 81788 60564 81844 62132
rect 82236 61684 82292 62636
rect 82348 62188 82404 63086
rect 82460 62578 82516 64204
rect 82460 62526 82462 62578
rect 82514 62526 82516 62578
rect 82460 62468 82516 62526
rect 82460 62402 82516 62412
rect 82348 62132 82516 62188
rect 82236 61590 82292 61628
rect 82348 60900 82404 60910
rect 82348 60806 82404 60844
rect 81452 60562 81844 60564
rect 81452 60510 81454 60562
rect 81506 60510 81844 60562
rect 81452 60508 81844 60510
rect 81900 60674 81956 60686
rect 81900 60622 81902 60674
rect 81954 60622 81956 60674
rect 81452 60452 81508 60508
rect 81452 60386 81508 60396
rect 81340 60162 81396 60172
rect 81676 60004 81732 60014
rect 81676 59910 81732 59948
rect 81116 59780 81172 59790
rect 81116 59444 81172 59724
rect 81900 59780 81956 60622
rect 82236 60564 82292 60574
rect 81900 59714 81956 59724
rect 82012 60004 82068 60014
rect 81276 59612 81540 59622
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81276 59546 81540 59556
rect 81228 59444 81284 59454
rect 81116 59442 81284 59444
rect 81116 59390 81230 59442
rect 81282 59390 81284 59442
rect 81116 59388 81284 59390
rect 81228 59378 81284 59388
rect 80220 58548 80276 58558
rect 81004 58548 81060 58716
rect 81676 59106 81732 59118
rect 81676 59054 81678 59106
rect 81730 59054 81732 59106
rect 81116 58548 81172 58558
rect 81004 58546 81172 58548
rect 81004 58494 81118 58546
rect 81170 58494 81172 58546
rect 81004 58492 81172 58494
rect 80220 58454 80276 58492
rect 81116 58482 81172 58492
rect 81564 58324 81620 58334
rect 81564 58230 81620 58268
rect 80668 58210 80724 58222
rect 80668 58158 80670 58210
rect 80722 58158 80724 58210
rect 80668 57988 80724 58158
rect 81676 58212 81732 59054
rect 82012 58436 82068 59948
rect 82124 59556 82180 59566
rect 82124 59442 82180 59500
rect 82124 59390 82126 59442
rect 82178 59390 82180 59442
rect 82124 58996 82180 59390
rect 82236 59108 82292 60508
rect 82460 60228 82516 62132
rect 82236 59042 82292 59052
rect 82348 60172 82516 60228
rect 82124 58930 82180 58940
rect 82012 58380 82292 58436
rect 81676 58146 81732 58156
rect 82124 58210 82180 58222
rect 82124 58158 82126 58210
rect 82178 58158 82180 58210
rect 81276 58044 81540 58054
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81276 57978 81540 57988
rect 80668 57922 80724 57932
rect 80332 57876 80388 57886
rect 80332 57762 80388 57820
rect 82012 57876 82068 57886
rect 82012 57782 82068 57820
rect 80332 57710 80334 57762
rect 80386 57710 80388 57762
rect 80332 57698 80388 57710
rect 80444 57764 80500 57774
rect 80668 57764 80724 57774
rect 80444 57762 80612 57764
rect 80444 57710 80446 57762
rect 80498 57710 80612 57762
rect 80444 57708 80612 57710
rect 80444 57698 80500 57708
rect 79996 56194 80052 57036
rect 80556 56980 80612 57708
rect 80668 57670 80724 57708
rect 81340 57764 81396 57774
rect 81340 57670 81396 57708
rect 81452 57764 81508 57774
rect 81452 57762 81620 57764
rect 81452 57710 81454 57762
rect 81506 57710 81620 57762
rect 81452 57708 81620 57710
rect 81452 57698 81508 57708
rect 81452 57426 81508 57438
rect 81452 57374 81454 57426
rect 81506 57374 81508 57426
rect 80556 56914 80612 56924
rect 81116 56980 81172 56990
rect 81116 56886 81172 56924
rect 80556 56644 80612 56654
rect 80332 56308 80388 56318
rect 80332 56214 80388 56252
rect 79996 56142 79998 56194
rect 80050 56142 80052 56194
rect 79996 56130 80052 56142
rect 79772 55916 80164 55972
rect 79772 55300 79828 55310
rect 79772 55206 79828 55244
rect 79996 51492 80052 51502
rect 79996 51398 80052 51436
rect 79884 51380 79940 51390
rect 79884 51286 79940 51324
rect 79996 51154 80052 51166
rect 79996 51102 79998 51154
rect 80050 51102 80052 51154
rect 79996 50428 80052 51102
rect 79212 49634 79268 49644
rect 79324 50372 79716 50428
rect 79772 50372 80052 50428
rect 79100 49028 79156 49038
rect 79100 48934 79156 48972
rect 78764 48302 78766 48354
rect 78818 48302 78820 48354
rect 78204 47348 78260 47358
rect 78764 47348 78820 48302
rect 78204 47346 78820 47348
rect 78204 47294 78206 47346
rect 78258 47294 78820 47346
rect 78204 47292 78820 47294
rect 78204 47282 78260 47292
rect 77980 46846 77982 46898
rect 78034 46846 78036 46898
rect 77980 46834 78036 46846
rect 79100 45780 79156 45790
rect 79100 45686 79156 45724
rect 78764 45668 78820 45678
rect 77756 45108 77812 45118
rect 77756 45014 77812 45052
rect 77420 44494 77422 44546
rect 77474 44494 77476 44546
rect 77420 44482 77476 44494
rect 77756 44436 77812 44446
rect 77756 44342 77812 44380
rect 77868 44212 77924 45612
rect 78428 45666 78820 45668
rect 78428 45614 78766 45666
rect 78818 45614 78820 45666
rect 78428 45612 78820 45614
rect 78428 45218 78484 45612
rect 78764 45602 78820 45612
rect 79212 45668 79268 45678
rect 78428 45166 78430 45218
rect 78482 45166 78484 45218
rect 78428 45154 78484 45166
rect 77980 44212 78036 44222
rect 77868 44210 78036 44212
rect 77868 44158 77982 44210
rect 78034 44158 78036 44210
rect 77868 44156 78036 44158
rect 77980 44146 78036 44156
rect 78540 44212 78596 44222
rect 78540 44118 78596 44156
rect 77756 43764 77812 43774
rect 77420 42980 77476 42990
rect 77420 42886 77476 42924
rect 77756 42978 77812 43708
rect 77868 43652 77924 43662
rect 77868 43558 77924 43596
rect 77756 42926 77758 42978
rect 77810 42926 77812 42978
rect 77756 42914 77812 42926
rect 79212 42866 79268 45612
rect 79324 43708 79380 50372
rect 79772 49138 79828 50372
rect 79772 49086 79774 49138
rect 79826 49086 79828 49138
rect 79772 49074 79828 49086
rect 80108 48468 80164 55916
rect 80556 55410 80612 56588
rect 81452 56644 81508 57374
rect 81564 56866 81620 57708
rect 81564 56814 81566 56866
rect 81618 56814 81620 56866
rect 81564 56802 81620 56814
rect 81788 56756 81844 56766
rect 81788 56662 81844 56700
rect 81900 56754 81956 56766
rect 81900 56702 81902 56754
rect 81954 56702 81956 56754
rect 81452 56578 81508 56588
rect 81900 56644 81956 56702
rect 81276 56476 81540 56486
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81276 56410 81540 56420
rect 81900 56308 81956 56588
rect 81900 56242 81956 56252
rect 80556 55358 80558 55410
rect 80610 55358 80612 55410
rect 80556 55346 80612 55358
rect 81788 55300 81844 55310
rect 81276 54908 81540 54918
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81276 54842 81540 54852
rect 80668 54516 80724 54526
rect 80556 54404 80612 54414
rect 80556 54310 80612 54348
rect 80220 53842 80276 53854
rect 80220 53790 80222 53842
rect 80274 53790 80276 53842
rect 80220 53172 80276 53790
rect 80220 53106 80276 53116
rect 80668 53508 80724 54460
rect 81788 54514 81844 55244
rect 82124 55300 82180 58158
rect 82124 55234 82180 55244
rect 81788 54462 81790 54514
rect 81842 54462 81844 54514
rect 81788 54450 81844 54462
rect 81340 54402 81396 54414
rect 81340 54350 81342 54402
rect 81394 54350 81396 54402
rect 81340 53508 81396 54350
rect 80668 53506 81396 53508
rect 80668 53454 80670 53506
rect 80722 53454 81396 53506
rect 80668 53452 81396 53454
rect 80556 51266 80612 51278
rect 80556 51214 80558 51266
rect 80610 51214 80612 51266
rect 80556 50148 80612 51214
rect 80668 50706 80724 53452
rect 81276 53340 81540 53350
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81276 53274 81540 53284
rect 81276 51772 81540 51782
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81276 51706 81540 51716
rect 82236 51604 82292 58380
rect 82348 56756 82404 60172
rect 82572 60116 82628 67116
rect 82796 66050 82852 66062
rect 82796 65998 82798 66050
rect 82850 65998 82852 66050
rect 82796 65716 82852 65998
rect 82796 65650 82852 65660
rect 82684 65378 82740 65390
rect 82684 65326 82686 65378
rect 82738 65326 82740 65378
rect 82684 65156 82740 65326
rect 82684 65090 82740 65100
rect 82908 65044 82964 69020
rect 83020 68628 83076 68638
rect 83020 67844 83076 68572
rect 83020 67750 83076 67788
rect 83132 67060 83188 69244
rect 83244 69234 83300 69244
rect 83356 69298 83412 70476
rect 83580 69412 83636 74508
rect 83804 74002 83860 75180
rect 83804 73950 83806 74002
rect 83858 73950 83860 74002
rect 83692 70754 83748 70766
rect 83692 70702 83694 70754
rect 83746 70702 83748 70754
rect 83692 70532 83748 70702
rect 83692 70466 83748 70476
rect 83580 69356 83748 69412
rect 83356 69246 83358 69298
rect 83410 69246 83412 69298
rect 83356 69234 83412 69246
rect 83580 69188 83636 69198
rect 83580 69094 83636 69132
rect 83468 68964 83524 68974
rect 83468 68514 83524 68908
rect 83468 68462 83470 68514
rect 83522 68462 83524 68514
rect 83244 67172 83300 67182
rect 83244 67078 83300 67116
rect 83132 66966 83188 67004
rect 83244 66834 83300 66846
rect 83244 66782 83246 66834
rect 83298 66782 83300 66834
rect 83244 66164 83300 66782
rect 83244 66098 83300 66108
rect 83244 65492 83300 65502
rect 83468 65492 83524 68462
rect 83692 67844 83748 69356
rect 83580 67730 83636 67742
rect 83580 67678 83582 67730
rect 83634 67678 83636 67730
rect 83580 67060 83636 67678
rect 83580 66994 83636 67004
rect 83692 67730 83748 67788
rect 83692 67678 83694 67730
rect 83746 67678 83748 67730
rect 83580 66052 83636 66062
rect 83580 65958 83636 65996
rect 83244 65490 83524 65492
rect 83244 65438 83246 65490
rect 83298 65438 83524 65490
rect 83244 65436 83524 65438
rect 83244 65426 83300 65436
rect 82908 64978 82964 64988
rect 83020 65268 83076 65278
rect 82684 64708 82740 64718
rect 82684 62692 82740 64652
rect 82908 64484 82964 64494
rect 82796 64482 82964 64484
rect 82796 64430 82910 64482
rect 82962 64430 82964 64482
rect 82796 64428 82964 64430
rect 82796 64372 82852 64428
rect 82908 64418 82964 64428
rect 82796 63924 82852 64316
rect 82908 64148 82964 64158
rect 82908 64054 82964 64092
rect 83020 64146 83076 65212
rect 83580 64932 83636 64942
rect 83020 64094 83022 64146
rect 83074 64094 83076 64146
rect 83020 64082 83076 64094
rect 83132 64820 83188 64830
rect 83132 64146 83188 64764
rect 83244 64708 83300 64718
rect 83244 64614 83300 64652
rect 83132 64094 83134 64146
rect 83186 64094 83188 64146
rect 83132 64082 83188 64094
rect 82796 63858 82852 63868
rect 83244 63922 83300 63934
rect 83244 63870 83246 63922
rect 83298 63870 83300 63922
rect 82908 63812 82964 63822
rect 82684 62626 82740 62636
rect 82796 63700 82852 63710
rect 82796 62466 82852 63644
rect 82796 62414 82798 62466
rect 82850 62414 82852 62466
rect 82796 62132 82852 62414
rect 82796 62066 82852 62076
rect 82684 61794 82740 61806
rect 82684 61742 82686 61794
rect 82738 61742 82740 61794
rect 82684 61682 82740 61742
rect 82684 61630 82686 61682
rect 82738 61630 82740 61682
rect 82684 61618 82740 61630
rect 82796 60900 82852 60910
rect 82796 60806 82852 60844
rect 82572 60060 82852 60116
rect 82460 60002 82516 60014
rect 82460 59950 82462 60002
rect 82514 59950 82516 60002
rect 82460 58994 82516 59950
rect 82572 59108 82628 59118
rect 82572 59014 82628 59052
rect 82460 58942 82462 58994
rect 82514 58942 82516 58994
rect 82460 58930 82516 58942
rect 82796 57764 82852 60060
rect 82348 56690 82404 56700
rect 82460 57708 82852 57764
rect 82348 53506 82404 53518
rect 82348 53454 82350 53506
rect 82402 53454 82404 53506
rect 82348 52500 82404 53454
rect 82348 52434 82404 52444
rect 82460 52276 82516 57708
rect 82908 57652 82964 63756
rect 83132 63700 83188 63710
rect 83020 63140 83076 63150
rect 83020 63046 83076 63084
rect 83020 62916 83076 62926
rect 83020 59444 83076 62860
rect 83132 61794 83188 63644
rect 83244 62580 83300 63870
rect 83244 62514 83300 62524
rect 83468 63922 83524 63934
rect 83468 63870 83470 63922
rect 83522 63870 83524 63922
rect 83244 62356 83300 62366
rect 83244 62262 83300 62300
rect 83468 62244 83524 63870
rect 83580 63924 83636 64876
rect 83580 63858 83636 63868
rect 83580 63026 83636 63038
rect 83580 62974 83582 63026
rect 83634 62974 83636 63026
rect 83580 62468 83636 62974
rect 83692 62804 83748 67678
rect 83804 67282 83860 73950
rect 84028 74900 84084 74910
rect 83916 72546 83972 72558
rect 83916 72494 83918 72546
rect 83970 72494 83972 72546
rect 83916 72324 83972 72494
rect 83916 68628 83972 72268
rect 83916 68562 83972 68572
rect 83804 67230 83806 67282
rect 83858 67230 83860 67282
rect 83804 67172 83860 67230
rect 83916 67618 83972 67630
rect 83916 67566 83918 67618
rect 83970 67566 83972 67618
rect 83916 67284 83972 67566
rect 83916 67218 83972 67228
rect 83804 67106 83860 67116
rect 84028 66388 84084 74844
rect 84252 74228 84308 75518
rect 84588 75682 84644 75694
rect 84588 75630 84590 75682
rect 84642 75630 84644 75682
rect 84588 75572 84644 75630
rect 84588 75506 84644 75516
rect 85260 75684 85316 75694
rect 85260 75570 85316 75628
rect 85260 75518 85262 75570
rect 85314 75518 85316 75570
rect 84364 75460 84420 75470
rect 84364 75458 84532 75460
rect 84364 75406 84366 75458
rect 84418 75406 84532 75458
rect 84364 75404 84532 75406
rect 84364 75394 84420 75404
rect 84476 74788 84532 75404
rect 85148 75124 85204 75134
rect 85260 75124 85316 75518
rect 85372 75570 85428 76300
rect 85596 75682 85652 77308
rect 85708 76692 85764 78766
rect 85932 78820 85988 81116
rect 86044 81106 86100 81116
rect 86492 80610 86548 80622
rect 86492 80558 86494 80610
rect 86546 80558 86548 80610
rect 86044 80500 86100 80510
rect 86044 80406 86100 80444
rect 86492 80498 86548 80558
rect 86492 80446 86494 80498
rect 86546 80446 86548 80498
rect 86492 80434 86548 80446
rect 86268 79716 86324 79726
rect 86268 79622 86324 79660
rect 86044 79604 86100 79614
rect 86044 79510 86100 79548
rect 85932 78754 85988 78764
rect 86156 78818 86212 78830
rect 86156 78766 86158 78818
rect 86210 78766 86212 78818
rect 86156 77252 86212 78766
rect 85708 76626 85764 76636
rect 86044 76916 86100 76926
rect 85596 75630 85598 75682
rect 85650 75630 85652 75682
rect 85596 75618 85652 75630
rect 86044 75796 86100 76860
rect 86044 75682 86100 75740
rect 86044 75630 86046 75682
rect 86098 75630 86100 75682
rect 86044 75618 86100 75630
rect 85372 75518 85374 75570
rect 85426 75518 85428 75570
rect 85372 75506 85428 75518
rect 86156 75570 86212 77196
rect 86156 75518 86158 75570
rect 86210 75518 86212 75570
rect 86156 75506 86212 75518
rect 86268 78594 86324 78606
rect 86268 78542 86270 78594
rect 86322 78542 86324 78594
rect 85148 75122 85316 75124
rect 85148 75070 85150 75122
rect 85202 75070 85316 75122
rect 85148 75068 85316 75070
rect 85148 75058 85204 75068
rect 84700 74788 84756 74798
rect 84476 74786 84756 74788
rect 84476 74734 84702 74786
rect 84754 74734 84756 74786
rect 84476 74732 84756 74734
rect 84700 74722 84756 74732
rect 84364 74228 84420 74238
rect 84252 74226 84420 74228
rect 84252 74174 84366 74226
rect 84418 74174 84420 74226
rect 84252 74172 84420 74174
rect 84364 74162 84420 74172
rect 84476 72324 84532 72334
rect 84476 72230 84532 72268
rect 85372 71876 85428 71886
rect 84252 71650 84308 71662
rect 84252 71598 84254 71650
rect 84306 71598 84308 71650
rect 84252 71204 84308 71598
rect 84252 71138 84308 71148
rect 85372 71202 85428 71820
rect 85372 71150 85374 71202
rect 85426 71150 85428 71202
rect 85372 71138 85428 71150
rect 85708 71204 85764 71214
rect 85708 71110 85764 71148
rect 86268 71092 86324 78542
rect 86380 76356 86436 76366
rect 86604 76356 86660 81228
rect 86716 80724 86772 81902
rect 86716 80658 86772 80668
rect 86828 81170 86884 82460
rect 86828 81118 86830 81170
rect 86882 81118 86884 81170
rect 86828 80500 86884 81118
rect 87388 80948 87444 83692
rect 87500 81170 87556 85148
rect 87724 84420 87780 84430
rect 87724 84326 87780 84364
rect 87612 83300 87668 83310
rect 87612 83206 87668 83244
rect 87500 81118 87502 81170
rect 87554 81118 87556 81170
rect 87500 81106 87556 81118
rect 87612 82628 87668 82638
rect 87612 81842 87668 82572
rect 87612 81790 87614 81842
rect 87666 81790 87668 81842
rect 87388 80892 87556 80948
rect 86828 79828 86884 80444
rect 86828 79604 86884 79772
rect 86716 79602 86884 79604
rect 86716 79550 86830 79602
rect 86882 79550 86884 79602
rect 86716 79548 86884 79550
rect 86716 78818 86772 79548
rect 86828 79538 86884 79548
rect 87388 79716 87444 79726
rect 86716 78766 86718 78818
rect 86770 78766 86772 78818
rect 86716 77140 86772 78766
rect 87388 77364 87444 79660
rect 87500 79602 87556 80892
rect 87500 79550 87502 79602
rect 87554 79550 87556 79602
rect 87500 79538 87556 79550
rect 87612 78988 87668 81790
rect 87612 78932 87780 78988
rect 87500 78820 87556 78830
rect 87500 78726 87556 78764
rect 87612 78036 87668 78046
rect 87612 77942 87668 77980
rect 87388 77308 87556 77364
rect 86716 77074 86772 77084
rect 87388 77138 87444 77150
rect 87388 77086 87390 77138
rect 87442 77086 87444 77138
rect 87276 76692 87332 76702
rect 87388 76692 87444 77086
rect 87276 76690 87444 76692
rect 87276 76638 87278 76690
rect 87330 76638 87444 76690
rect 87276 76636 87444 76638
rect 87276 76626 87332 76636
rect 87052 76578 87108 76590
rect 87052 76526 87054 76578
rect 87106 76526 87108 76578
rect 86940 76466 86996 76478
rect 86940 76414 86942 76466
rect 86994 76414 86996 76466
rect 86604 76300 86884 76356
rect 86380 76262 86436 76300
rect 86716 75796 86772 75806
rect 86716 75702 86772 75740
rect 86380 75684 86436 75694
rect 86380 75590 86436 75628
rect 86604 72548 86660 72558
rect 86604 72322 86660 72492
rect 86604 72270 86606 72322
rect 86658 72270 86660 72322
rect 86268 71036 86436 71092
rect 85932 70868 85988 70878
rect 85932 70774 85988 70812
rect 86268 70866 86324 70878
rect 86268 70814 86270 70866
rect 86322 70814 86324 70866
rect 84588 70756 84644 70766
rect 84588 70662 84644 70700
rect 85372 70084 85428 70094
rect 85372 69990 85428 70028
rect 85596 70084 85652 70094
rect 84364 69634 84420 69646
rect 84364 69582 84366 69634
rect 84418 69582 84420 69634
rect 84364 69524 84420 69582
rect 84364 69458 84420 69468
rect 84476 69412 84532 69422
rect 84476 69318 84532 69356
rect 85260 69410 85316 69422
rect 85260 69358 85262 69410
rect 85314 69358 85316 69410
rect 84364 69188 84420 69198
rect 84364 69094 84420 69132
rect 85260 68964 85316 69358
rect 84252 67844 84308 67854
rect 84252 67750 84308 67788
rect 85260 67842 85316 68908
rect 85260 67790 85262 67842
rect 85314 67790 85316 67842
rect 85260 67778 85316 67790
rect 85148 67732 85204 67742
rect 84252 67396 84308 67406
rect 84252 67170 84308 67340
rect 84252 67118 84254 67170
rect 84306 67118 84308 67170
rect 84252 67106 84308 67118
rect 84700 67396 84756 67406
rect 84700 67170 84756 67340
rect 84700 67118 84702 67170
rect 84754 67118 84756 67170
rect 84700 67106 84756 67118
rect 85148 67170 85204 67676
rect 85148 67118 85150 67170
rect 85202 67118 85204 67170
rect 85148 67106 85204 67118
rect 85260 67620 85316 67630
rect 85148 66388 85204 66398
rect 85260 66388 85316 67564
rect 85372 67284 85428 67294
rect 85372 67190 85428 67228
rect 85484 67172 85540 67182
rect 85484 67078 85540 67116
rect 84028 66322 84084 66332
rect 84476 66386 85316 66388
rect 84476 66334 85150 66386
rect 85202 66334 85316 66386
rect 84476 66332 85316 66334
rect 84252 66164 84308 66174
rect 84252 66070 84308 66108
rect 84364 66162 84420 66174
rect 84364 66110 84366 66162
rect 84418 66110 84420 66162
rect 84028 66050 84084 66062
rect 84028 65998 84030 66050
rect 84082 65998 84084 66050
rect 83916 65492 83972 65502
rect 84028 65492 84084 65998
rect 83916 65490 84084 65492
rect 83916 65438 83918 65490
rect 83970 65438 84084 65490
rect 83916 65436 84084 65438
rect 84140 66052 84196 66062
rect 84140 65604 84196 65996
rect 84364 65716 84420 66110
rect 84364 65650 84420 65660
rect 83916 65426 83972 65436
rect 84140 64594 84196 65548
rect 84476 65044 84532 66332
rect 85148 66322 85204 66332
rect 84252 64988 84532 65044
rect 85372 66276 85428 66286
rect 85372 65828 85428 66220
rect 84252 64706 84308 64988
rect 85372 64708 85428 65772
rect 84252 64654 84254 64706
rect 84306 64654 84308 64706
rect 84252 64642 84308 64654
rect 85036 64652 85428 64708
rect 84140 64542 84142 64594
rect 84194 64542 84196 64594
rect 84140 64530 84196 64542
rect 83916 64484 83972 64494
rect 83916 64482 84084 64484
rect 83916 64430 83918 64482
rect 83970 64430 84084 64482
rect 83916 64428 84084 64430
rect 83916 64418 83972 64428
rect 83916 63924 83972 63934
rect 83916 63830 83972 63868
rect 83804 63028 83860 63038
rect 83804 62934 83860 62972
rect 83916 62916 83972 62926
rect 83916 62822 83972 62860
rect 83692 62748 83860 62804
rect 83580 62402 83636 62412
rect 83692 62356 83748 62366
rect 83692 62262 83748 62300
rect 83468 62178 83524 62188
rect 83804 61908 83860 62748
rect 84028 62468 84084 64428
rect 85036 64146 85092 64652
rect 85372 64594 85428 64652
rect 85484 66052 85540 66062
rect 85484 64706 85540 65996
rect 85484 64654 85486 64706
rect 85538 64654 85540 64706
rect 85484 64642 85540 64654
rect 85372 64542 85374 64594
rect 85426 64542 85428 64594
rect 85372 64530 85428 64542
rect 85148 64484 85204 64494
rect 85484 64484 85540 64494
rect 85148 64482 85316 64484
rect 85148 64430 85150 64482
rect 85202 64430 85316 64482
rect 85148 64428 85316 64430
rect 85148 64418 85204 64428
rect 85036 64094 85038 64146
rect 85090 64094 85092 64146
rect 85036 64082 85092 64094
rect 84812 64036 84868 64046
rect 84812 63942 84868 63980
rect 84924 63924 84980 63934
rect 85148 63924 85204 63934
rect 84980 63868 85092 63924
rect 84924 63858 84980 63868
rect 84364 63810 84420 63822
rect 84364 63758 84366 63810
rect 84418 63758 84420 63810
rect 84364 63252 84420 63758
rect 84364 63186 84420 63196
rect 84028 62402 84084 62412
rect 84252 63138 84308 63150
rect 84252 63086 84254 63138
rect 84306 63086 84308 63138
rect 83132 61742 83134 61794
rect 83186 61742 83188 61794
rect 83132 61730 83188 61742
rect 83580 61852 83860 61908
rect 83916 62356 83972 62366
rect 83468 61572 83524 61582
rect 83468 61478 83524 61516
rect 83244 60788 83300 60798
rect 83244 60694 83300 60732
rect 83580 60564 83636 61852
rect 83692 61684 83748 61694
rect 83692 61570 83748 61628
rect 83804 61684 83860 61694
rect 83916 61684 83972 62300
rect 83804 61682 83972 61684
rect 83804 61630 83806 61682
rect 83858 61630 83972 61682
rect 83804 61628 83972 61630
rect 83804 61618 83860 61628
rect 83692 61518 83694 61570
rect 83746 61518 83748 61570
rect 83692 61506 83748 61518
rect 83916 61460 83972 61470
rect 83804 61458 83972 61460
rect 83804 61406 83918 61458
rect 83970 61406 83972 61458
rect 83804 61404 83972 61406
rect 83580 60508 83748 60564
rect 83580 60340 83636 60350
rect 83132 60116 83188 60126
rect 83132 60022 83188 60060
rect 83580 60114 83636 60284
rect 83580 60062 83582 60114
rect 83634 60062 83636 60114
rect 83580 60050 83636 60062
rect 83132 59444 83188 59454
rect 83020 59442 83188 59444
rect 83020 59390 83134 59442
rect 83186 59390 83188 59442
rect 83020 59388 83188 59390
rect 83132 59378 83188 59388
rect 83468 59444 83524 59454
rect 83132 58660 83188 58670
rect 83132 58546 83188 58604
rect 83132 58494 83134 58546
rect 83186 58494 83188 58546
rect 83132 58482 83188 58494
rect 83468 58658 83524 59388
rect 83468 58606 83470 58658
rect 83522 58606 83524 58658
rect 83468 58548 83524 58606
rect 83580 58548 83636 58558
rect 83468 58546 83636 58548
rect 83468 58494 83582 58546
rect 83634 58494 83636 58546
rect 83468 58492 83636 58494
rect 83580 58482 83636 58492
rect 83692 57764 83748 60508
rect 83580 57708 83748 57764
rect 83804 57764 83860 61404
rect 83916 61394 83972 61404
rect 84252 61124 84308 63086
rect 84476 63028 84532 63038
rect 84364 62580 84420 62590
rect 84364 62486 84420 62524
rect 84364 61348 84420 61358
rect 84364 61254 84420 61292
rect 84252 61058 84308 61068
rect 84140 60900 84196 60910
rect 84028 60844 84140 60900
rect 84028 60340 84084 60844
rect 84140 60768 84196 60844
rect 84252 60788 84308 60798
rect 84252 60694 84308 60732
rect 84140 60564 84196 60574
rect 84476 60564 84532 62972
rect 84700 62580 84756 62590
rect 84588 62466 84644 62478
rect 84588 62414 84590 62466
rect 84642 62414 84644 62466
rect 84588 61348 84644 62414
rect 84588 60900 84644 61292
rect 84588 60834 84644 60844
rect 84700 62354 84756 62524
rect 85036 62468 85092 63868
rect 85148 63830 85204 63868
rect 85260 63140 85316 64428
rect 85260 63074 85316 63084
rect 85372 63812 85428 63822
rect 85148 62916 85204 62926
rect 85372 62916 85428 63756
rect 85148 62914 85428 62916
rect 85148 62862 85150 62914
rect 85202 62862 85428 62914
rect 85148 62860 85428 62862
rect 85148 62692 85204 62860
rect 85148 62626 85204 62636
rect 85148 62468 85204 62478
rect 85036 62466 85204 62468
rect 85036 62414 85150 62466
rect 85202 62414 85204 62466
rect 85036 62412 85204 62414
rect 85148 62402 85204 62412
rect 84700 62302 84702 62354
rect 84754 62302 84756 62354
rect 84140 60562 84532 60564
rect 84140 60510 84142 60562
rect 84194 60510 84532 60562
rect 84140 60508 84532 60510
rect 84140 60498 84196 60508
rect 84084 60284 84196 60340
rect 84028 60274 84084 60284
rect 83916 60228 83972 60238
rect 83916 60116 83972 60172
rect 84028 60116 84084 60126
rect 83916 60114 84084 60116
rect 83916 60062 84030 60114
rect 84082 60062 84084 60114
rect 83916 60060 84084 60062
rect 84028 60050 84084 60060
rect 82908 57650 83188 57652
rect 82908 57598 82910 57650
rect 82962 57598 83188 57650
rect 82908 57596 83188 57598
rect 82908 57586 82964 57596
rect 82572 57540 82628 57550
rect 82572 57538 82852 57540
rect 82572 57486 82574 57538
rect 82626 57486 82852 57538
rect 82572 57484 82852 57486
rect 82572 57474 82628 57484
rect 82684 56756 82740 56766
rect 82572 56642 82628 56654
rect 82572 56590 82574 56642
rect 82626 56590 82628 56642
rect 82572 55412 82628 56590
rect 82572 55346 82628 55356
rect 82684 55410 82740 56700
rect 82796 56644 82852 57484
rect 82796 56578 82852 56588
rect 82908 57316 82964 57326
rect 82684 55358 82686 55410
rect 82738 55358 82740 55410
rect 82684 55346 82740 55358
rect 82796 56084 82852 56094
rect 82572 54628 82628 54638
rect 82572 54534 82628 54572
rect 82684 52388 82740 52398
rect 82460 52220 82628 52276
rect 82460 51604 82516 51614
rect 82236 51602 82516 51604
rect 82236 51550 82462 51602
rect 82514 51550 82516 51602
rect 82236 51548 82516 51550
rect 81228 51492 81284 51502
rect 81228 51398 81284 51436
rect 81452 51492 81508 51502
rect 81452 51398 81508 51436
rect 81900 51492 81956 51502
rect 80668 50654 80670 50706
rect 80722 50654 80724 50706
rect 80668 50642 80724 50654
rect 81564 51378 81620 51390
rect 81564 51326 81566 51378
rect 81618 51326 81620 51378
rect 81564 51156 81620 51326
rect 81564 50372 81620 51100
rect 81564 50306 81620 50316
rect 81676 50484 81732 50494
rect 81276 50204 81540 50214
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81276 50138 81540 50148
rect 80444 49700 80500 49710
rect 80444 49606 80500 49644
rect 80556 49588 80612 50092
rect 81676 50036 81732 50428
rect 80556 49522 80612 49532
rect 81340 49980 81732 50036
rect 81340 49698 81396 49980
rect 81340 49646 81342 49698
rect 81394 49646 81396 49698
rect 81340 48804 81396 49646
rect 81788 49810 81844 49822
rect 81788 49758 81790 49810
rect 81842 49758 81844 49810
rect 80108 48402 80164 48412
rect 81116 48748 81396 48804
rect 81676 49028 81732 49038
rect 79548 48242 79604 48254
rect 79548 48190 79550 48242
rect 79602 48190 79604 48242
rect 79324 43652 79492 43708
rect 79212 42814 79214 42866
rect 79266 42814 79268 42866
rect 79212 42802 79268 42814
rect 77756 42756 77812 42766
rect 77756 42194 77812 42700
rect 77980 42756 78036 42766
rect 77980 42642 78036 42700
rect 77980 42590 77982 42642
rect 78034 42590 78036 42642
rect 77980 42578 78036 42590
rect 78540 42644 78596 42654
rect 78540 42550 78596 42588
rect 77756 42142 77758 42194
rect 77810 42142 77812 42194
rect 77756 42084 77812 42142
rect 77308 42028 77476 42084
rect 76860 41916 77140 41972
rect 76860 41858 76916 41916
rect 76860 41806 76862 41858
rect 76914 41806 76916 41858
rect 76860 41748 76916 41806
rect 77308 41858 77364 41870
rect 77308 41806 77310 41858
rect 77362 41806 77364 41858
rect 77308 41748 77364 41806
rect 77420 41860 77476 42028
rect 77756 42018 77812 42028
rect 77420 41794 77476 41804
rect 78204 41860 78260 41870
rect 76860 41692 77140 41748
rect 76636 41580 77028 41636
rect 76524 41300 76580 41310
rect 76300 40964 76356 40974
rect 76300 40870 76356 40908
rect 76412 39620 76468 39630
rect 76412 39526 76468 39564
rect 76188 38948 76244 38958
rect 76188 38854 76244 38892
rect 76524 38162 76580 41244
rect 76524 38110 76526 38162
rect 76578 38110 76580 38162
rect 76524 38052 76580 38110
rect 76524 37986 76580 37996
rect 76076 36482 76132 36540
rect 76076 36430 76078 36482
rect 76130 36430 76132 36482
rect 76076 36418 76132 36430
rect 76412 37378 76468 37390
rect 76412 37326 76414 37378
rect 76466 37326 76468 37378
rect 76412 36932 76468 37326
rect 76412 36370 76468 36876
rect 76412 36318 76414 36370
rect 76466 36318 76468 36370
rect 74956 36260 75012 36270
rect 74732 35924 74788 35934
rect 74732 35698 74788 35868
rect 74956 35810 75012 36204
rect 76412 36260 76468 36318
rect 76412 36194 76468 36204
rect 74956 35758 74958 35810
rect 75010 35758 75012 35810
rect 74956 35746 75012 35758
rect 75292 35924 75348 35934
rect 74732 35646 74734 35698
rect 74786 35646 74788 35698
rect 74732 35634 74788 35646
rect 75292 34354 75348 35868
rect 76524 35812 76580 35822
rect 76524 35718 76580 35756
rect 76748 35698 76804 35710
rect 76748 35646 76750 35698
rect 76802 35646 76804 35698
rect 75852 35588 75908 35598
rect 76748 35588 76804 35646
rect 75852 35586 76804 35588
rect 75852 35534 75854 35586
rect 75906 35534 76804 35586
rect 75852 35532 76804 35534
rect 75852 35522 75908 35532
rect 75516 35474 75572 35486
rect 75516 35422 75518 35474
rect 75570 35422 75572 35474
rect 75516 35028 75572 35422
rect 75516 34962 75572 34972
rect 76524 35028 76580 35038
rect 76524 34934 76580 34972
rect 75292 34302 75294 34354
rect 75346 34302 75348 34354
rect 75292 34290 75348 34302
rect 74620 34130 75124 34132
rect 74620 34078 74622 34130
rect 74674 34078 75124 34130
rect 74620 34076 75124 34078
rect 74620 34066 74676 34076
rect 73724 32788 73780 33292
rect 73836 33852 74452 33908
rect 73836 33124 73892 33852
rect 74284 33346 74340 33358
rect 74284 33294 74286 33346
rect 74338 33294 74340 33346
rect 74284 33236 74340 33294
rect 74732 33348 74788 33358
rect 74732 33254 74788 33292
rect 74284 33170 74340 33180
rect 73836 33058 73892 33068
rect 73836 32788 73892 32798
rect 73724 32732 73836 32788
rect 73836 32656 73892 32732
rect 74284 32788 74340 32798
rect 74284 32694 74340 32732
rect 75068 32786 75124 34076
rect 75964 34018 76020 34030
rect 75964 33966 75966 34018
rect 76018 33966 76020 34018
rect 75740 33122 75796 33134
rect 75740 33070 75742 33122
rect 75794 33070 75796 33122
rect 75068 32734 75070 32786
rect 75122 32734 75124 32786
rect 75068 32722 75124 32734
rect 75516 32788 75572 32798
rect 75740 32788 75796 33070
rect 75572 32732 75796 32788
rect 75516 32694 75572 32732
rect 75964 32676 76020 33966
rect 76300 33348 76356 33358
rect 76188 32676 76244 32686
rect 75964 32620 76188 32676
rect 76188 32582 76244 32620
rect 73500 31892 73780 31948
rect 73724 31890 73780 31892
rect 73724 31838 73726 31890
rect 73778 31838 73780 31890
rect 73724 31826 73780 31838
rect 76300 31892 76356 33292
rect 76748 32788 76804 32798
rect 76748 32694 76804 32732
rect 76412 31892 76468 31902
rect 76300 31890 76468 31892
rect 76300 31838 76414 31890
rect 76466 31838 76468 31890
rect 76300 31836 76468 31838
rect 76412 31826 76468 31836
rect 76972 25284 77028 41580
rect 77084 37940 77140 41692
rect 77308 41300 77364 41692
rect 77308 41244 77476 41300
rect 77308 41076 77364 41086
rect 77308 40982 77364 41020
rect 77196 40404 77252 40414
rect 77196 39730 77252 40348
rect 77196 39678 77198 39730
rect 77250 39678 77252 39730
rect 77196 39666 77252 39678
rect 77084 37490 77140 37884
rect 77084 37438 77086 37490
rect 77138 37438 77140 37490
rect 77084 37426 77140 37438
rect 77308 39620 77364 39630
rect 77308 38050 77364 39564
rect 77308 37998 77310 38050
rect 77362 37998 77364 38050
rect 77308 37156 77364 37998
rect 77420 37492 77476 41244
rect 77532 41186 77588 41198
rect 77532 41134 77534 41186
rect 77586 41134 77588 41186
rect 77532 38836 77588 41134
rect 77532 38770 77588 38780
rect 77756 40516 77812 40526
rect 77756 40290 77812 40460
rect 78204 40516 78260 41804
rect 78204 40450 78260 40460
rect 78988 41074 79044 41086
rect 78988 41022 78990 41074
rect 79042 41022 79044 41074
rect 77756 40238 77758 40290
rect 77810 40238 77812 40290
rect 77756 39396 77812 40238
rect 78428 39618 78484 39630
rect 78428 39566 78430 39618
rect 78482 39566 78484 39618
rect 77868 39396 77924 39406
rect 78428 39396 78484 39566
rect 77756 39394 78484 39396
rect 77756 39342 77870 39394
rect 77922 39342 78484 39394
rect 77756 39340 78484 39342
rect 77756 38164 77812 39340
rect 77868 39330 77924 39340
rect 78988 39058 79044 41022
rect 79324 40962 79380 40974
rect 79324 40910 79326 40962
rect 79378 40910 79380 40962
rect 79212 39732 79268 39742
rect 79324 39732 79380 40910
rect 79212 39730 79380 39732
rect 79212 39678 79214 39730
rect 79266 39678 79380 39730
rect 79212 39676 79380 39678
rect 79212 39666 79268 39676
rect 78988 39006 78990 39058
rect 79042 39006 79044 39058
rect 78988 38994 79044 39006
rect 78316 38724 78372 38734
rect 78316 38630 78372 38668
rect 79324 38724 79380 38734
rect 79324 38630 79380 38668
rect 77420 37436 77588 37492
rect 77420 37156 77476 37166
rect 77308 37154 77476 37156
rect 77308 37102 77422 37154
rect 77474 37102 77476 37154
rect 77308 37100 77476 37102
rect 77420 37090 77476 37100
rect 77196 36932 77252 36942
rect 77196 36596 77252 36876
rect 77532 36932 77588 37436
rect 77532 36866 77588 36876
rect 77420 36596 77476 36606
rect 77196 36594 77364 36596
rect 77196 36542 77198 36594
rect 77250 36542 77364 36594
rect 77196 36540 77364 36542
rect 77196 36530 77252 36540
rect 77308 35922 77364 36540
rect 77308 35870 77310 35922
rect 77362 35870 77364 35922
rect 77308 35858 77364 35870
rect 77084 35028 77140 35038
rect 77084 32562 77140 34972
rect 77308 34916 77364 34926
rect 77308 34822 77364 34860
rect 77308 33234 77364 33246
rect 77308 33182 77310 33234
rect 77362 33182 77364 33234
rect 77308 32788 77364 33182
rect 77308 32722 77364 32732
rect 77084 32510 77086 32562
rect 77138 32510 77140 32562
rect 77084 32498 77140 32510
rect 77420 31948 77476 36540
rect 77644 36596 77700 36606
rect 77644 36502 77700 36540
rect 77756 34916 77812 38108
rect 78988 38164 79044 38174
rect 78988 38070 79044 38108
rect 77868 38052 77924 38062
rect 77868 37958 77924 37996
rect 78540 38052 78596 38062
rect 78540 37958 78596 37996
rect 77868 37380 77924 37390
rect 77868 37286 77924 37324
rect 77756 34850 77812 34860
rect 78764 34914 78820 34926
rect 78764 34862 78766 34914
rect 78818 34862 78820 34914
rect 77532 34356 77588 34366
rect 77532 33348 77588 34300
rect 78764 34132 78820 34862
rect 78092 34020 78148 34030
rect 77532 32562 77588 33292
rect 77644 34018 78148 34020
rect 77644 33966 78094 34018
rect 78146 33966 78148 34018
rect 77644 33964 78148 33966
rect 77644 33234 77700 33964
rect 78092 33954 78148 33964
rect 77644 33182 77646 33234
rect 77698 33182 77700 33234
rect 77644 33170 77700 33182
rect 77868 33572 77924 33582
rect 77532 32510 77534 32562
rect 77586 32510 77588 32562
rect 77868 32676 77924 33516
rect 78316 33348 78372 33358
rect 78764 33348 78820 34076
rect 79436 33684 79492 43652
rect 79548 43428 79604 48190
rect 80444 48242 80500 48254
rect 80444 48190 80446 48242
rect 80498 48190 80500 48242
rect 80444 44996 80500 48190
rect 81004 47572 81060 47582
rect 81004 47478 81060 47516
rect 81004 46564 81060 46574
rect 80668 45780 80724 45790
rect 80668 45686 80724 45724
rect 80668 45108 80724 45118
rect 80556 44996 80612 45006
rect 80444 44994 80612 44996
rect 80444 44942 80558 44994
rect 80610 44942 80612 44994
rect 80444 44940 80612 44942
rect 80444 44212 80500 44940
rect 80556 44930 80612 44940
rect 80668 44434 80724 45052
rect 80668 44382 80670 44434
rect 80722 44382 80724 44434
rect 80668 44370 80724 44382
rect 80444 44146 80500 44156
rect 79996 43428 80052 43438
rect 79548 43426 80052 43428
rect 79548 43374 79998 43426
rect 80050 43374 80052 43426
rect 79548 43372 80052 43374
rect 79548 42644 79604 43372
rect 79996 43362 80052 43372
rect 79548 42578 79604 42588
rect 80556 42868 80612 42878
rect 80556 41300 80612 42812
rect 80556 41234 80612 41244
rect 80444 40404 80500 40414
rect 80444 40310 80500 40348
rect 80108 38948 80164 38958
rect 80108 38854 80164 38892
rect 79996 38834 80052 38846
rect 79996 38782 79998 38834
rect 80050 38782 80052 38834
rect 79996 38052 80052 38782
rect 79996 37828 80052 37996
rect 79996 37762 80052 37772
rect 79548 34802 79604 34814
rect 79548 34750 79550 34802
rect 79602 34750 79604 34802
rect 79548 34354 79604 34750
rect 79548 34302 79550 34354
rect 79602 34302 79604 34354
rect 79548 34290 79604 34302
rect 79884 34244 79940 34254
rect 79884 34150 79940 34188
rect 79436 33618 79492 33628
rect 78316 33346 78820 33348
rect 78316 33294 78318 33346
rect 78370 33294 78820 33346
rect 78316 33292 78820 33294
rect 80668 33348 80724 33358
rect 78316 33282 78372 33292
rect 78988 33234 79044 33246
rect 78988 33182 78990 33234
rect 79042 33182 79044 33234
rect 78988 32788 79044 33182
rect 78988 32722 79044 32732
rect 80668 32786 80724 33292
rect 80668 32734 80670 32786
rect 80722 32734 80724 32786
rect 80668 32722 80724 32734
rect 77868 32544 77924 32620
rect 77532 32498 77588 32510
rect 81004 31948 81060 46508
rect 81116 45332 81172 48748
rect 81276 48636 81540 48646
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81276 48570 81540 48580
rect 81676 48242 81732 48972
rect 81676 48190 81678 48242
rect 81730 48190 81732 48242
rect 81676 47572 81732 48190
rect 81788 47684 81844 49758
rect 81900 49138 81956 51436
rect 82236 51492 82292 51548
rect 82460 51538 82516 51548
rect 82236 51426 82292 51436
rect 82012 51266 82068 51278
rect 82012 51214 82014 51266
rect 82066 51214 82068 51266
rect 82012 51156 82068 51214
rect 82012 51090 82068 51100
rect 82348 50148 82404 50158
rect 82348 50034 82404 50092
rect 82348 49982 82350 50034
rect 82402 49982 82404 50034
rect 82348 49970 82404 49982
rect 82236 49812 82292 49822
rect 82236 49718 82292 49756
rect 81900 49086 81902 49138
rect 81954 49086 81956 49138
rect 81900 49074 81956 49086
rect 82348 48804 82404 48814
rect 81788 47618 81844 47628
rect 82236 48802 82404 48804
rect 82236 48750 82350 48802
rect 82402 48750 82404 48802
rect 82236 48748 82404 48750
rect 81676 47506 81732 47516
rect 82236 47572 82292 48748
rect 82348 48738 82404 48748
rect 82348 48356 82404 48366
rect 82348 48262 82404 48300
rect 82236 47478 82292 47516
rect 81276 47068 81540 47078
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81276 47002 81540 47012
rect 82460 46900 82516 46910
rect 82572 46900 82628 52220
rect 82460 46898 82572 46900
rect 82460 46846 82462 46898
rect 82514 46846 82572 46898
rect 82460 46844 82572 46846
rect 82460 46834 82516 46844
rect 82572 46768 82628 46844
rect 82236 46674 82292 46686
rect 82236 46622 82238 46674
rect 82290 46622 82292 46674
rect 81676 46564 81732 46574
rect 81676 46470 81732 46508
rect 82236 46564 82292 46622
rect 82236 46498 82292 46508
rect 81340 45892 81396 45902
rect 82236 45892 82292 45902
rect 81340 45890 82292 45892
rect 81340 45838 81342 45890
rect 81394 45838 82238 45890
rect 82290 45838 82292 45890
rect 81340 45836 82292 45838
rect 81340 45826 81396 45836
rect 82236 45826 82292 45836
rect 82572 45892 82628 45902
rect 82572 45798 82628 45836
rect 82684 45780 82740 52332
rect 82796 50596 82852 56028
rect 82796 50530 82852 50540
rect 82796 48802 82852 48814
rect 82796 48750 82798 48802
rect 82850 48750 82852 48802
rect 82796 48356 82852 48750
rect 82796 48290 82852 48300
rect 82796 45780 82852 45790
rect 82684 45724 82796 45780
rect 81564 45668 81620 45678
rect 81564 45666 82180 45668
rect 81564 45614 81566 45666
rect 81618 45614 82180 45666
rect 82796 45648 82852 45724
rect 81564 45612 82180 45614
rect 81564 45602 81620 45612
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 81116 45276 81732 45332
rect 81116 45108 81172 45118
rect 81116 41972 81172 45052
rect 81340 45108 81396 45118
rect 81340 45014 81396 45052
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 81340 41972 81396 41982
rect 81116 41970 81396 41972
rect 81116 41918 81342 41970
rect 81394 41918 81396 41970
rect 81116 41916 81396 41918
rect 81340 41906 81396 41916
rect 81564 41076 81620 41086
rect 81564 40982 81620 41020
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 81228 40404 81284 40414
rect 81228 40310 81284 40348
rect 81340 39732 81396 39742
rect 81116 39676 81340 39732
rect 81116 39060 81172 39676
rect 81340 39638 81396 39676
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 81340 39060 81396 39070
rect 81116 39058 81396 39060
rect 81116 39006 81342 39058
rect 81394 39006 81396 39058
rect 81116 39004 81396 39006
rect 81116 38948 81172 39004
rect 81340 38994 81396 39004
rect 81452 39060 81508 39070
rect 81116 38882 81172 38892
rect 81452 38050 81508 39004
rect 81452 37998 81454 38050
rect 81506 37998 81508 38050
rect 81452 37986 81508 37998
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 81228 35924 81284 35934
rect 81228 35830 81284 35868
rect 81676 35922 81732 45276
rect 82124 45218 82180 45612
rect 82124 45166 82126 45218
rect 82178 45166 82180 45218
rect 82124 45154 82180 45166
rect 81788 42756 81844 42766
rect 81788 42754 81956 42756
rect 81788 42702 81790 42754
rect 81842 42702 81956 42754
rect 81788 42700 81956 42702
rect 81788 42690 81844 42700
rect 81900 41860 81956 42700
rect 82012 42530 82068 42542
rect 82012 42478 82014 42530
rect 82066 42478 82068 42530
rect 82012 42084 82068 42478
rect 82124 42084 82180 42094
rect 82012 42082 82180 42084
rect 82012 42030 82126 42082
rect 82178 42030 82180 42082
rect 82012 42028 82180 42030
rect 82124 42018 82180 42028
rect 81900 41804 82180 41860
rect 82124 41410 82180 41804
rect 82124 41358 82126 41410
rect 82178 41358 82180 41410
rect 82124 41346 82180 41358
rect 82460 41186 82516 41198
rect 82460 41134 82462 41186
rect 82514 41134 82516 41186
rect 81676 35870 81678 35922
rect 81730 35870 81732 35922
rect 81676 35026 81732 35870
rect 81788 41076 81844 41086
rect 81788 36820 81844 41020
rect 82460 40292 82516 41134
rect 82684 41076 82740 41086
rect 82684 40982 82740 41020
rect 82460 40226 82516 40236
rect 82684 40402 82740 40414
rect 82684 40350 82686 40402
rect 82738 40350 82740 40402
rect 82684 40180 82740 40350
rect 82348 39620 82404 39630
rect 82684 39620 82740 40124
rect 82908 39732 82964 57260
rect 83132 56868 83188 57596
rect 83468 57428 83524 57438
rect 83244 56868 83300 56878
rect 83132 56866 83300 56868
rect 83132 56814 83246 56866
rect 83298 56814 83300 56866
rect 83132 56812 83300 56814
rect 83020 56644 83076 56654
rect 83020 54852 83076 56588
rect 83244 55748 83300 56812
rect 83468 56754 83524 57372
rect 83468 56702 83470 56754
rect 83522 56702 83524 56754
rect 83468 56690 83524 56702
rect 83244 55682 83300 55692
rect 83356 55412 83412 55422
rect 83020 54786 83076 54796
rect 83132 55300 83188 55310
rect 83020 53620 83076 53630
rect 83020 53526 83076 53564
rect 83020 53172 83076 53182
rect 83132 53172 83188 55244
rect 83356 55298 83412 55356
rect 83356 55246 83358 55298
rect 83410 55246 83412 55298
rect 83356 53844 83412 55246
rect 83356 53778 83412 53788
rect 83580 55186 83636 57708
rect 83804 57698 83860 57708
rect 83916 59106 83972 59118
rect 83916 59054 83918 59106
rect 83970 59054 83972 59106
rect 83916 58994 83972 59054
rect 83916 58942 83918 58994
rect 83970 58942 83972 58994
rect 83692 57540 83748 57550
rect 83692 57538 83860 57540
rect 83692 57486 83694 57538
rect 83746 57486 83860 57538
rect 83692 57484 83860 57486
rect 83692 57474 83748 57484
rect 83580 55134 83582 55186
rect 83634 55134 83636 55186
rect 83020 53170 83188 53172
rect 83020 53118 83022 53170
rect 83074 53118 83188 53170
rect 83020 53116 83188 53118
rect 83244 53730 83300 53742
rect 83244 53678 83246 53730
rect 83298 53678 83300 53730
rect 83020 53106 83076 53116
rect 83244 52388 83300 53678
rect 83580 53620 83636 55134
rect 83804 57204 83860 57484
rect 83916 57316 83972 58942
rect 84028 58660 84084 58670
rect 84028 57650 84084 58604
rect 84140 58546 84196 60284
rect 84364 60004 84420 60014
rect 84364 59442 84420 59948
rect 84476 59892 84532 59902
rect 84476 59798 84532 59836
rect 84364 59390 84366 59442
rect 84418 59390 84420 59442
rect 84364 59378 84420 59390
rect 84140 58494 84142 58546
rect 84194 58494 84196 58546
rect 84140 58482 84196 58494
rect 84476 59108 84532 59118
rect 84476 58658 84532 59052
rect 84476 58606 84478 58658
rect 84530 58606 84532 58658
rect 84476 58546 84532 58606
rect 84476 58494 84478 58546
rect 84530 58494 84532 58546
rect 84476 58482 84532 58494
rect 84028 57598 84030 57650
rect 84082 57598 84084 57650
rect 84028 57586 84084 57598
rect 84476 57988 84532 57998
rect 84700 57988 84756 62302
rect 85484 61684 85540 64428
rect 85260 61572 85316 61582
rect 85260 61478 85316 61516
rect 85484 61570 85540 61628
rect 85484 61518 85486 61570
rect 85538 61518 85540 61570
rect 85484 61506 85540 61518
rect 85596 61012 85652 70028
rect 86268 70084 86324 70814
rect 86268 70018 86324 70028
rect 86380 69860 86436 71036
rect 86380 69794 86436 69804
rect 85708 69748 85764 69758
rect 85708 62580 85764 69692
rect 86044 69524 86100 69534
rect 86044 69430 86100 69468
rect 85820 68852 85876 68862
rect 85820 67396 85876 68796
rect 86044 67732 86100 67742
rect 86044 67638 86100 67676
rect 85820 67060 85876 67340
rect 86492 67284 86548 67322
rect 86492 67218 86548 67228
rect 86380 67060 86436 67070
rect 85820 67058 86436 67060
rect 85820 67006 86382 67058
rect 86434 67006 86436 67058
rect 85820 67004 86436 67006
rect 85820 66274 85876 67004
rect 86380 66994 86436 67004
rect 85820 66222 85822 66274
rect 85874 66222 85876 66274
rect 85820 66210 85876 66222
rect 85932 66052 85988 66062
rect 85932 66050 86100 66052
rect 85932 65998 85934 66050
rect 85986 65998 86100 66050
rect 85932 65996 86100 65998
rect 85932 65986 85988 65996
rect 86044 65378 86100 65996
rect 86156 66050 86212 66062
rect 86156 65998 86158 66050
rect 86210 65998 86212 66050
rect 86156 65716 86212 65998
rect 86492 66052 86548 66062
rect 86492 65958 86548 65996
rect 86156 65650 86212 65660
rect 86044 65326 86046 65378
rect 86098 65326 86100 65378
rect 86044 65314 86100 65326
rect 86604 64820 86660 72270
rect 86716 67172 86772 67182
rect 86716 67078 86772 67116
rect 86828 66948 86884 76300
rect 86940 75684 86996 76414
rect 86940 75618 86996 75628
rect 87052 75572 87108 76526
rect 87052 75506 87108 75516
rect 87164 72548 87220 72558
rect 87164 72454 87220 72492
rect 87052 70754 87108 70766
rect 87052 70702 87054 70754
rect 87106 70702 87108 70754
rect 87052 70084 87108 70702
rect 87164 70196 87220 70206
rect 87164 70102 87220 70140
rect 87052 70018 87108 70028
rect 87164 69860 87220 69870
rect 87052 66948 87108 66958
rect 86828 66946 87108 66948
rect 86828 66894 87054 66946
rect 87106 66894 87108 66946
rect 86828 66892 87108 66894
rect 86716 65604 86772 65614
rect 86716 65510 86772 65548
rect 86828 65602 86884 66892
rect 87052 66882 87108 66892
rect 86828 65550 86830 65602
rect 86882 65550 86884 65602
rect 86828 65538 86884 65550
rect 87052 66276 87108 66286
rect 86716 65268 86772 65278
rect 86716 65174 86772 65212
rect 86604 64764 86772 64820
rect 86044 64594 86100 64606
rect 86044 64542 86046 64594
rect 86098 64542 86100 64594
rect 85932 63924 85988 63934
rect 85820 63026 85876 63038
rect 85820 62974 85822 63026
rect 85874 62974 85876 63026
rect 85820 62916 85876 62974
rect 85820 62850 85876 62860
rect 85932 62692 85988 63868
rect 86044 63922 86100 64542
rect 86044 63870 86046 63922
rect 86098 63870 86100 63922
rect 86044 63812 86100 63870
rect 86268 64594 86324 64606
rect 86268 64542 86270 64594
rect 86322 64542 86324 64594
rect 86268 64148 86324 64542
rect 86604 64594 86660 64606
rect 86604 64542 86606 64594
rect 86658 64542 86660 64594
rect 86268 63924 86324 64092
rect 86268 63792 86324 63868
rect 86380 64482 86436 64494
rect 86380 64430 86382 64482
rect 86434 64430 86436 64482
rect 86044 63746 86100 63756
rect 86156 63252 86212 63262
rect 86156 63158 86212 63196
rect 86268 63140 86324 63150
rect 86268 63046 86324 63084
rect 86044 63028 86100 63038
rect 86044 62934 86100 62972
rect 85932 62636 86324 62692
rect 85708 62524 86212 62580
rect 86044 62356 86100 62366
rect 86156 62356 86212 62524
rect 86268 62578 86324 62636
rect 86268 62526 86270 62578
rect 86322 62526 86324 62578
rect 86268 62514 86324 62526
rect 86380 62580 86436 64430
rect 86604 64148 86660 64542
rect 86604 64082 86660 64092
rect 86604 63922 86660 63934
rect 86604 63870 86606 63922
rect 86658 63870 86660 63922
rect 86492 63810 86548 63822
rect 86492 63758 86494 63810
rect 86546 63758 86548 63810
rect 86492 63138 86548 63758
rect 86492 63086 86494 63138
rect 86546 63086 86548 63138
rect 86492 63074 86548 63086
rect 86604 63028 86660 63870
rect 86604 62962 86660 62972
rect 86604 62580 86660 62590
rect 86380 62578 86660 62580
rect 86380 62526 86606 62578
rect 86658 62526 86660 62578
rect 86380 62524 86660 62526
rect 86604 62514 86660 62524
rect 86380 62356 86436 62366
rect 86156 62354 86436 62356
rect 86156 62302 86382 62354
rect 86434 62302 86436 62354
rect 86156 62300 86436 62302
rect 86044 62262 86100 62300
rect 86380 62290 86436 62300
rect 86492 62356 86548 62366
rect 86492 62262 86548 62300
rect 85708 62244 85764 62254
rect 85708 61682 85764 62188
rect 85708 61630 85710 61682
rect 85762 61630 85764 61682
rect 85708 61618 85764 61630
rect 86268 61796 86324 61806
rect 86268 61682 86324 61740
rect 86268 61630 86270 61682
rect 86322 61630 86324 61682
rect 86268 61618 86324 61630
rect 85932 61572 85988 61582
rect 86716 61572 86772 64764
rect 87052 64818 87108 66220
rect 87164 66052 87220 69804
rect 87388 68628 87444 68638
rect 87388 68534 87444 68572
rect 87500 67620 87556 77308
rect 87612 76692 87668 76702
rect 87724 76692 87780 78876
rect 87612 76690 87780 76692
rect 87612 76638 87614 76690
rect 87666 76638 87780 76690
rect 87612 76636 87780 76638
rect 87612 76626 87668 76636
rect 87836 74116 87892 74126
rect 87724 70980 87780 70990
rect 87836 70980 87892 74060
rect 88060 73220 88116 85708
rect 89180 85764 89236 86380
rect 89292 86434 89348 86446
rect 89292 86382 89294 86434
rect 89346 86382 89348 86434
rect 89292 86324 89348 86382
rect 89292 86258 89348 86268
rect 89180 85762 89348 85764
rect 89180 85710 89182 85762
rect 89234 85710 89348 85762
rect 89180 85708 89348 85710
rect 89180 85698 89236 85708
rect 88844 85316 88900 85326
rect 88844 85222 88900 85260
rect 88172 85204 88228 85214
rect 88172 85110 88228 85148
rect 89180 85204 89236 85214
rect 89180 85110 89236 85148
rect 89292 85092 89348 85708
rect 89628 85092 89684 85102
rect 89292 85090 89684 85092
rect 89292 85038 89630 85090
rect 89682 85038 89684 85090
rect 89292 85036 89684 85038
rect 89292 84420 89348 84430
rect 89292 84326 89348 84364
rect 88508 84308 88564 84318
rect 88284 84084 88340 84094
rect 88284 83746 88340 84028
rect 88284 83694 88286 83746
rect 88338 83694 88340 83746
rect 88284 83682 88340 83694
rect 88396 83524 88452 83534
rect 88396 81170 88452 83468
rect 88396 81118 88398 81170
rect 88450 81118 88452 81170
rect 88396 81106 88452 81118
rect 88508 80500 88564 84252
rect 89516 84306 89572 84318
rect 89516 84254 89518 84306
rect 89570 84254 89572 84306
rect 89404 84196 89460 84206
rect 88620 83748 88676 83758
rect 88620 83654 88676 83692
rect 88844 83410 88900 83422
rect 88844 83358 88846 83410
rect 88898 83358 88900 83410
rect 88844 83300 88900 83358
rect 89404 83410 89460 84140
rect 89516 84084 89572 84254
rect 89516 84018 89572 84028
rect 89404 83358 89406 83410
rect 89458 83358 89460 83410
rect 89404 83346 89460 83358
rect 88844 83234 88900 83244
rect 89628 83300 89684 85036
rect 89740 84978 89796 86492
rect 91196 86546 91588 86548
rect 91196 86494 91534 86546
rect 91586 86494 91588 86546
rect 91196 86492 91588 86494
rect 89740 84926 89742 84978
rect 89794 84926 89796 84978
rect 89740 84914 89796 84926
rect 90636 85762 90692 85774
rect 90636 85710 90638 85762
rect 90690 85710 90692 85762
rect 90524 84868 90580 84878
rect 90412 84866 90580 84868
rect 90412 84814 90526 84866
rect 90578 84814 90580 84866
rect 90412 84812 90580 84814
rect 90188 84308 90244 84318
rect 90188 84214 90244 84252
rect 89628 83234 89684 83244
rect 90412 82628 90468 84812
rect 90524 84802 90580 84812
rect 90524 84532 90580 84542
rect 90524 83634 90580 84476
rect 90636 84196 90692 85710
rect 91196 85314 91252 86492
rect 91532 86482 91588 86492
rect 91868 86546 91924 88844
rect 93772 88898 93828 88910
rect 93772 88846 93774 88898
rect 93826 88846 93828 88898
rect 91868 86494 91870 86546
rect 91922 86494 91924 86546
rect 91868 86482 91924 86494
rect 92652 87444 92708 87454
rect 91196 85262 91198 85314
rect 91250 85262 91252 85314
rect 91196 85250 91252 85262
rect 91532 86324 91588 86334
rect 91196 85092 91252 85102
rect 90636 84140 90804 84196
rect 90524 83582 90526 83634
rect 90578 83582 90580 83634
rect 90524 83570 90580 83582
rect 90748 83524 90804 84140
rect 90748 83458 90804 83468
rect 90972 84194 91028 84206
rect 90972 84142 90974 84194
rect 91026 84142 91028 84194
rect 90972 83188 91028 84142
rect 91196 83746 91252 85036
rect 91532 85092 91588 86268
rect 91532 85090 91700 85092
rect 91532 85038 91534 85090
rect 91586 85038 91700 85090
rect 91532 85036 91700 85038
rect 91532 85026 91588 85036
rect 91532 84196 91588 84206
rect 91532 84102 91588 84140
rect 91196 83694 91198 83746
rect 91250 83694 91252 83746
rect 91196 83682 91252 83694
rect 91532 83524 91588 83534
rect 91532 83430 91588 83468
rect 91644 83188 91700 85036
rect 92204 85090 92260 85102
rect 92204 85038 92206 85090
rect 92258 85038 92260 85090
rect 92204 84532 92260 85038
rect 92204 83524 92260 84476
rect 92204 83430 92260 83468
rect 92316 84980 92372 84990
rect 92316 83410 92372 84924
rect 92316 83358 92318 83410
rect 92370 83358 92372 83410
rect 92316 83346 92372 83358
rect 90972 83132 92036 83188
rect 90412 82562 90468 82572
rect 90636 82626 90692 82638
rect 90636 82574 90638 82626
rect 90690 82574 90692 82626
rect 90636 82348 90692 82574
rect 90636 82292 90804 82348
rect 90748 81732 90804 82292
rect 90972 81732 91028 81742
rect 90748 81730 91028 81732
rect 90748 81678 90974 81730
rect 91026 81678 91028 81730
rect 90748 81676 91028 81678
rect 90972 80724 91028 81676
rect 90972 80658 91028 80668
rect 91196 80724 91252 80734
rect 88508 80498 88900 80500
rect 88508 80446 88510 80498
rect 88562 80446 88900 80498
rect 88508 80444 88900 80446
rect 88508 80434 88564 80444
rect 88396 79940 88452 79950
rect 88396 79602 88452 79884
rect 88396 79550 88398 79602
rect 88450 79550 88452 79602
rect 88396 79538 88452 79550
rect 88844 78932 88900 80444
rect 89628 79940 89684 79950
rect 89180 79828 89236 79838
rect 89180 79734 89236 79772
rect 89628 79826 89684 79884
rect 89628 79774 89630 79826
rect 89682 79774 89684 79826
rect 89628 79762 89684 79774
rect 90412 79490 90468 79502
rect 90412 79438 90414 79490
rect 90466 79438 90468 79490
rect 88956 78932 89012 78942
rect 88844 78930 89012 78932
rect 88844 78878 88958 78930
rect 89010 78878 89012 78930
rect 88844 78876 89012 78878
rect 88396 78818 88452 78830
rect 88396 78766 88398 78818
rect 88450 78766 88452 78818
rect 88396 78596 88452 78766
rect 88396 78530 88452 78540
rect 88396 78036 88452 78046
rect 88844 78036 88900 78876
rect 88956 78866 89012 78876
rect 90412 78820 90468 79438
rect 90412 78754 90468 78764
rect 89516 78596 89572 78606
rect 89516 78502 89572 78540
rect 89404 78146 89460 78158
rect 89404 78094 89406 78146
rect 89458 78094 89460 78146
rect 88172 78034 88900 78036
rect 88172 77982 88398 78034
rect 88450 77982 88900 78034
rect 88172 77980 88900 77982
rect 89180 78036 89236 78046
rect 88172 77250 88228 77980
rect 88396 77970 88452 77980
rect 88732 77362 88788 77980
rect 89180 77942 89236 77980
rect 88732 77310 88734 77362
rect 88786 77310 88788 77362
rect 88732 77298 88788 77310
rect 89404 77364 89460 78094
rect 89516 78148 89572 78158
rect 89516 78054 89572 78092
rect 89404 77298 89460 77308
rect 88172 77198 88174 77250
rect 88226 77198 88228 77250
rect 88172 77186 88228 77198
rect 90860 77026 90916 77038
rect 90860 76974 90862 77026
rect 90914 76974 90916 77026
rect 90300 76578 90356 76590
rect 90300 76526 90302 76578
rect 90354 76526 90356 76578
rect 90300 75794 90356 76526
rect 90300 75742 90302 75794
rect 90354 75742 90356 75794
rect 90300 75730 90356 75742
rect 90636 76466 90692 76478
rect 90636 76414 90638 76466
rect 90690 76414 90692 76466
rect 89516 75682 89572 75694
rect 89516 75630 89518 75682
rect 89570 75630 89572 75682
rect 89068 75458 89124 75470
rect 89068 75406 89070 75458
rect 89122 75406 89124 75458
rect 88508 75010 88564 75022
rect 88508 74958 88510 75010
rect 88562 74958 88564 75010
rect 88284 74900 88340 74910
rect 88284 74806 88340 74844
rect 88508 74228 88564 74958
rect 89068 74676 89124 75406
rect 89404 74900 89460 74910
rect 89404 74806 89460 74844
rect 89068 74610 89124 74620
rect 88620 74228 88676 74238
rect 88508 74226 88676 74228
rect 88508 74174 88622 74226
rect 88674 74174 88676 74226
rect 88508 74172 88676 74174
rect 88620 74162 88676 74172
rect 89516 74116 89572 75630
rect 90636 75236 90692 76414
rect 90860 76468 90916 76974
rect 91196 76468 91252 80668
rect 91420 79716 91476 79726
rect 91420 77922 91476 79660
rect 91868 79492 91924 79502
rect 91644 79380 91700 79390
rect 91644 78818 91700 79324
rect 91644 78766 91646 78818
rect 91698 78766 91700 78818
rect 91644 78754 91700 78766
rect 91868 78706 91924 79436
rect 91980 78988 92036 83132
rect 92652 82740 92708 87388
rect 93548 85874 93604 85886
rect 93548 85822 93550 85874
rect 93602 85822 93604 85874
rect 92764 85764 92820 85774
rect 92764 85762 93268 85764
rect 92764 85710 92766 85762
rect 92818 85710 93268 85762
rect 92764 85708 93268 85710
rect 92764 85698 92820 85708
rect 93212 84978 93268 85708
rect 93548 85204 93604 85822
rect 93548 85138 93604 85148
rect 93436 85092 93492 85102
rect 93436 84998 93492 85036
rect 93212 84926 93214 84978
rect 93266 84926 93268 84978
rect 93212 84914 93268 84926
rect 93772 84980 93828 88846
rect 96636 88620 96900 88630
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96636 88554 96900 88564
rect 94556 87444 94612 87454
rect 94556 87350 94612 87388
rect 95116 87444 95172 87454
rect 95116 87350 95172 87388
rect 96636 87052 96900 87062
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96636 86986 96900 86996
rect 95564 86548 95620 86558
rect 95116 86546 95620 86548
rect 95116 86494 95566 86546
rect 95618 86494 95620 86546
rect 95116 86492 95620 86494
rect 93772 84914 93828 84924
rect 94892 85204 94948 85214
rect 94892 85090 94948 85148
rect 94892 85038 94894 85090
rect 94946 85038 94948 85090
rect 94444 84866 94500 84878
rect 94444 84814 94446 84866
rect 94498 84814 94500 84866
rect 94444 84532 94500 84814
rect 94108 84476 94444 84532
rect 93660 84194 93716 84206
rect 93660 84142 93662 84194
rect 93714 84142 93716 84194
rect 93324 83522 93380 83534
rect 93324 83470 93326 83522
rect 93378 83470 93380 83522
rect 92652 82738 93156 82740
rect 92652 82686 92654 82738
rect 92706 82686 93156 82738
rect 92652 82684 93156 82686
rect 92652 82674 92708 82684
rect 92428 81732 92484 81742
rect 92204 81676 92428 81732
rect 92204 81394 92260 81676
rect 92428 81638 92484 81676
rect 92204 81342 92206 81394
rect 92258 81342 92260 81394
rect 92204 81284 92260 81342
rect 92204 81218 92260 81228
rect 92876 80946 92932 80958
rect 92876 80894 92878 80946
rect 92930 80894 92932 80946
rect 92428 80724 92484 80734
rect 92428 80386 92484 80668
rect 92428 80334 92430 80386
rect 92482 80334 92484 80386
rect 92428 80322 92484 80334
rect 92540 79492 92596 79502
rect 92540 79398 92596 79436
rect 92876 78988 92932 80894
rect 93100 80724 93156 82684
rect 93324 82178 93380 83470
rect 93548 83412 93604 83422
rect 93660 83412 93716 84142
rect 93548 83410 93716 83412
rect 93548 83358 93550 83410
rect 93602 83358 93716 83410
rect 93548 83356 93716 83358
rect 93548 83346 93604 83356
rect 94108 82292 94164 84476
rect 94444 84466 94500 84476
rect 94444 84306 94500 84318
rect 94444 84254 94446 84306
rect 94498 84254 94500 84306
rect 93324 82126 93326 82178
rect 93378 82126 93380 82178
rect 93324 82114 93380 82126
rect 93772 82236 94164 82292
rect 93660 81956 93716 81966
rect 93772 81956 93828 82236
rect 94108 82068 94164 82236
rect 94108 82002 94164 82012
rect 94220 84196 94276 84206
rect 93660 81954 93828 81956
rect 93660 81902 93662 81954
rect 93714 81902 93828 81954
rect 93660 81900 93828 81902
rect 93548 81282 93604 81294
rect 93548 81230 93550 81282
rect 93602 81230 93604 81282
rect 93212 81060 93268 81070
rect 93212 80966 93268 81004
rect 93100 80498 93156 80668
rect 93100 80446 93102 80498
rect 93154 80446 93156 80498
rect 93100 80434 93156 80446
rect 93548 80724 93604 81230
rect 93548 80498 93604 80668
rect 93548 80446 93550 80498
rect 93602 80446 93604 80498
rect 93548 80434 93604 80446
rect 93324 80388 93380 80398
rect 93324 79602 93380 80332
rect 93324 79550 93326 79602
rect 93378 79550 93380 79602
rect 93324 79538 93380 79550
rect 93660 78988 93716 81900
rect 93884 81842 93940 81854
rect 93884 81790 93886 81842
rect 93938 81790 93940 81842
rect 93884 81732 93940 81790
rect 94220 81842 94276 84140
rect 94332 83636 94388 83646
rect 94332 83542 94388 83580
rect 94444 83524 94500 84254
rect 94892 83524 94948 85038
rect 94444 83522 94948 83524
rect 94444 83470 94894 83522
rect 94946 83470 94948 83522
rect 94444 83468 94948 83470
rect 94220 81790 94222 81842
rect 94274 81790 94276 81842
rect 94220 81778 94276 81790
rect 94892 82626 94948 83468
rect 94892 82574 94894 82626
rect 94946 82574 94948 82626
rect 93772 81282 93828 81294
rect 93772 81230 93774 81282
rect 93826 81230 93828 81282
rect 93772 79716 93828 81230
rect 93884 80724 93940 81676
rect 94668 81060 94724 81070
rect 94724 81004 94836 81060
rect 94668 80928 94724 81004
rect 93884 80658 93940 80668
rect 94556 80724 94612 80734
rect 94332 80276 94388 80286
rect 94388 80220 94500 80276
rect 94332 80182 94388 80220
rect 93772 79650 93828 79660
rect 93996 79380 94052 79390
rect 93996 79286 94052 79324
rect 94332 79378 94388 79390
rect 94332 79326 94334 79378
rect 94386 79326 94388 79378
rect 91980 78932 92148 78988
rect 92876 78932 93268 78988
rect 93660 78932 93828 78988
rect 91868 78654 91870 78706
rect 91922 78654 91924 78706
rect 91868 78642 91924 78654
rect 91420 77870 91422 77922
rect 91474 77870 91476 77922
rect 91420 77858 91476 77870
rect 91868 76468 91924 76478
rect 90860 76466 91924 76468
rect 90860 76414 91870 76466
rect 91922 76414 91924 76466
rect 90860 76412 91924 76414
rect 90636 75170 90692 75180
rect 91420 75236 91476 75246
rect 91420 75122 91476 75180
rect 91420 75070 91422 75122
rect 91474 75070 91476 75122
rect 91420 75058 91476 75070
rect 89964 75010 90020 75022
rect 89964 74958 89966 75010
rect 90018 74958 90020 75010
rect 89740 74788 89796 74798
rect 89740 74694 89796 74732
rect 89516 74050 89572 74060
rect 89964 74676 90020 74958
rect 89964 74228 90020 74620
rect 89740 74004 89796 74014
rect 88172 73444 88228 73454
rect 88172 73442 88452 73444
rect 88172 73390 88174 73442
rect 88226 73390 88452 73442
rect 88172 73388 88452 73390
rect 88172 73378 88228 73388
rect 88060 73164 88340 73220
rect 87724 70978 87892 70980
rect 87724 70926 87726 70978
rect 87778 70926 87892 70978
rect 87724 70924 87892 70926
rect 88060 70980 88116 70990
rect 87724 70914 87780 70924
rect 88060 70418 88116 70924
rect 88060 70366 88062 70418
rect 88114 70366 88116 70418
rect 88060 70354 88116 70366
rect 87724 70082 87780 70094
rect 87724 70030 87726 70082
rect 87778 70030 87780 70082
rect 87724 68852 87780 70030
rect 88172 69522 88228 69534
rect 88172 69470 88174 69522
rect 88226 69470 88228 69522
rect 88172 69300 88228 69470
rect 88172 69234 88228 69244
rect 87724 68786 87780 68796
rect 88284 68404 88340 73164
rect 88396 71090 88452 73388
rect 88508 73332 88564 73342
rect 88508 73238 88564 73276
rect 89404 73332 89460 73342
rect 89404 73238 89460 73276
rect 89740 73106 89796 73948
rect 89964 73442 90020 74172
rect 89964 73390 89966 73442
rect 90018 73390 90020 73442
rect 89964 73378 90020 73390
rect 90524 75010 90580 75022
rect 90524 74958 90526 75010
rect 90578 74958 90580 75010
rect 90524 74228 90580 74958
rect 90860 74788 90916 74798
rect 90748 74228 90804 74238
rect 90524 74226 90804 74228
rect 90524 74174 90750 74226
rect 90802 74174 90804 74226
rect 90524 74172 90804 74174
rect 90524 73442 90580 74172
rect 90748 74162 90804 74172
rect 90524 73390 90526 73442
rect 90578 73390 90580 73442
rect 90524 73378 90580 73390
rect 89740 73054 89742 73106
rect 89794 73054 89796 73106
rect 88396 71038 88398 71090
rect 88450 71038 88452 71090
rect 88396 71026 88452 71038
rect 89180 72434 89236 72446
rect 89180 72382 89182 72434
rect 89234 72382 89236 72434
rect 89180 71764 89236 72382
rect 89180 70644 89236 71708
rect 88956 70588 89236 70644
rect 89292 71204 89348 71214
rect 88508 70084 88564 70094
rect 88956 70084 89012 70588
rect 89292 70418 89348 71148
rect 89292 70366 89294 70418
rect 89346 70366 89348 70418
rect 89292 70354 89348 70366
rect 89404 70980 89460 70990
rect 89740 70980 89796 73054
rect 89852 71764 89908 71774
rect 89852 71670 89908 71708
rect 90860 71204 90916 74732
rect 91756 74676 91812 74686
rect 91532 74620 91756 74676
rect 91532 74340 91588 74620
rect 91756 74544 91812 74620
rect 91420 74284 91588 74340
rect 91084 74228 91140 74238
rect 91084 73554 91140 74172
rect 91308 74004 91364 74014
rect 91308 73910 91364 73948
rect 91084 73502 91086 73554
rect 91138 73502 91140 73554
rect 91084 73490 91140 73502
rect 90524 71090 90580 71102
rect 90524 71038 90526 71090
rect 90578 71038 90580 71090
rect 90524 70980 90580 71038
rect 89740 70924 90580 70980
rect 90860 70980 90916 71148
rect 88508 70082 89012 70084
rect 88508 70030 88510 70082
rect 88562 70030 89012 70082
rect 88508 70028 89012 70030
rect 88508 68628 88564 70028
rect 89068 69412 89124 69422
rect 89068 69318 89124 69356
rect 88732 69298 88788 69310
rect 88732 69246 88734 69298
rect 88786 69246 88788 69298
rect 88732 68852 88788 69246
rect 88844 69300 88900 69310
rect 88844 69206 88900 69244
rect 88732 68786 88788 68796
rect 88508 68562 88564 68572
rect 89404 68626 89460 70924
rect 89628 70196 89684 70272
rect 89684 70140 89796 70196
rect 89628 70130 89684 70140
rect 89628 69972 89684 69982
rect 89404 68574 89406 68626
rect 89458 68574 89460 68626
rect 89404 68562 89460 68574
rect 89516 69522 89572 69534
rect 89516 69470 89518 69522
rect 89570 69470 89572 69522
rect 89516 68740 89572 69470
rect 88284 68348 88900 68404
rect 87500 67554 87556 67564
rect 88172 67954 88228 67966
rect 88172 67902 88174 67954
rect 88226 67902 88228 67954
rect 88172 67284 88228 67902
rect 88172 67218 88228 67228
rect 88732 67954 88788 67966
rect 88732 67902 88734 67954
rect 88786 67902 88788 67954
rect 87724 67172 87780 67182
rect 87724 67078 87780 67116
rect 88732 67172 88788 67902
rect 88732 67106 88788 67116
rect 87836 67060 87892 67070
rect 87836 66966 87892 67004
rect 88284 66946 88340 66958
rect 88284 66894 88286 66946
rect 88338 66894 88340 66946
rect 87724 66836 87780 66846
rect 87724 66834 88116 66836
rect 87724 66782 87726 66834
rect 87778 66782 88116 66834
rect 87724 66780 88116 66782
rect 87724 66770 87780 66780
rect 88060 66386 88116 66780
rect 88060 66334 88062 66386
rect 88114 66334 88116 66386
rect 88060 66322 88116 66334
rect 87388 66276 87444 66286
rect 87388 66182 87444 66220
rect 87948 66276 88004 66286
rect 87164 65986 87220 65996
rect 87388 65380 87444 65390
rect 87388 65378 87780 65380
rect 87388 65326 87390 65378
rect 87442 65326 87780 65378
rect 87388 65324 87780 65326
rect 87388 65314 87444 65324
rect 87052 64766 87054 64818
rect 87106 64766 87108 64818
rect 87052 64146 87108 64766
rect 87500 64148 87556 64158
rect 87052 64094 87054 64146
rect 87106 64094 87108 64146
rect 87052 64082 87108 64094
rect 87276 64146 87556 64148
rect 87276 64094 87502 64146
rect 87554 64094 87556 64146
rect 87276 64092 87556 64094
rect 87276 63924 87332 64092
rect 87500 64082 87556 64092
rect 87612 64036 87668 64046
rect 87052 63868 87332 63924
rect 87388 63924 87444 63934
rect 87052 63700 87108 63868
rect 86940 62914 86996 62926
rect 86940 62862 86942 62914
rect 86994 62862 86996 62914
rect 86940 62804 86996 62862
rect 86940 62738 86996 62748
rect 85932 61570 86212 61572
rect 85932 61518 85934 61570
rect 85986 61518 86212 61570
rect 85932 61516 86212 61518
rect 85932 61506 85988 61516
rect 85484 60956 85652 61012
rect 85820 61124 85876 61134
rect 85820 61010 85876 61068
rect 85820 60958 85822 61010
rect 85874 60958 85876 61010
rect 85148 60786 85204 60798
rect 85148 60734 85150 60786
rect 85202 60734 85204 60786
rect 84812 60676 84868 60686
rect 84812 60674 84980 60676
rect 84812 60622 84814 60674
rect 84866 60622 84980 60674
rect 84812 60620 84980 60622
rect 84812 60610 84868 60620
rect 84812 60004 84868 60014
rect 84812 59106 84868 59948
rect 84812 59054 84814 59106
rect 84866 59054 84868 59106
rect 84812 58660 84868 59054
rect 84812 58594 84868 58604
rect 84924 58324 84980 60620
rect 85148 60116 85204 60734
rect 85148 58546 85204 60060
rect 85260 59892 85316 59902
rect 85260 59890 85428 59892
rect 85260 59838 85262 59890
rect 85314 59838 85428 59890
rect 85260 59836 85428 59838
rect 85260 59826 85316 59836
rect 85148 58494 85150 58546
rect 85202 58494 85204 58546
rect 85148 58482 85204 58494
rect 85260 59108 85316 59118
rect 84924 58258 84980 58268
rect 84476 57650 84532 57932
rect 84476 57598 84478 57650
rect 84530 57598 84532 57650
rect 84476 57586 84532 57598
rect 84588 57932 84756 57988
rect 83916 57250 83972 57260
rect 83804 55076 83860 57148
rect 84028 56866 84084 56878
rect 84028 56814 84030 56866
rect 84082 56814 84084 56866
rect 84028 56196 84084 56814
rect 84364 56644 84420 56654
rect 84364 56642 84532 56644
rect 84364 56590 84366 56642
rect 84418 56590 84532 56642
rect 84364 56588 84532 56590
rect 84364 56578 84420 56588
rect 83804 55010 83860 55020
rect 83916 56140 84084 56196
rect 83916 54404 83972 56140
rect 84028 55970 84084 55982
rect 84028 55918 84030 55970
rect 84082 55918 84084 55970
rect 84028 55300 84084 55918
rect 84364 55300 84420 55310
rect 84028 55234 84084 55244
rect 84252 55298 84420 55300
rect 84252 55246 84366 55298
rect 84418 55246 84420 55298
rect 84252 55244 84420 55246
rect 84140 55074 84196 55086
rect 84140 55022 84142 55074
rect 84194 55022 84196 55074
rect 84140 54628 84196 55022
rect 84140 54562 84196 54572
rect 83804 53956 83860 53966
rect 83916 53956 83972 54348
rect 83804 53954 83972 53956
rect 83804 53902 83806 53954
rect 83858 53902 83972 53954
rect 83804 53900 83972 53902
rect 84140 53956 84196 53966
rect 84252 53956 84308 55244
rect 84364 55234 84420 55244
rect 84140 53954 84308 53956
rect 84140 53902 84142 53954
rect 84194 53902 84308 53954
rect 84140 53900 84308 53902
rect 84364 55076 84420 55086
rect 83804 53890 83860 53900
rect 84140 53890 84196 53900
rect 83580 53554 83636 53564
rect 83244 52322 83300 52332
rect 83804 50596 83860 50606
rect 83804 50502 83860 50540
rect 84364 50428 84420 55020
rect 84476 54628 84532 56588
rect 84476 54562 84532 54572
rect 84364 50372 84532 50428
rect 83020 49810 83076 49822
rect 83020 49758 83022 49810
rect 83074 49758 83076 49810
rect 83020 49588 83076 49758
rect 83580 49810 83636 49822
rect 83580 49758 83582 49810
rect 83634 49758 83636 49810
rect 83580 49700 83636 49758
rect 83580 49634 83636 49644
rect 83804 49812 83860 49822
rect 83020 49522 83076 49532
rect 83132 48916 83188 48926
rect 83580 48916 83636 48926
rect 83132 48914 83636 48916
rect 83132 48862 83134 48914
rect 83186 48862 83582 48914
rect 83634 48862 83636 48914
rect 83132 48860 83636 48862
rect 83132 48850 83188 48860
rect 83580 48850 83636 48860
rect 83804 48916 83860 49756
rect 84364 49812 84420 49822
rect 84364 49718 84420 49756
rect 84140 49588 84196 49598
rect 83916 49476 83972 49486
rect 83916 49026 83972 49420
rect 83916 48974 83918 49026
rect 83970 48974 83972 49026
rect 83916 48962 83972 48974
rect 83020 48804 83076 48814
rect 83804 48784 83860 48860
rect 83020 47572 83076 48748
rect 83468 47572 83524 47582
rect 83020 47570 83524 47572
rect 83020 47518 83470 47570
rect 83522 47518 83524 47570
rect 83020 47516 83524 47518
rect 83468 47506 83524 47516
rect 84140 47570 84196 49532
rect 84364 49476 84420 49486
rect 84364 49138 84420 49420
rect 84364 49086 84366 49138
rect 84418 49086 84420 49138
rect 84364 49028 84420 49086
rect 84364 48962 84420 48972
rect 84476 48580 84532 50372
rect 84588 50148 84644 57932
rect 84700 57764 84756 57774
rect 84700 57670 84756 57708
rect 85260 57650 85316 59052
rect 85372 58548 85428 59836
rect 85372 58482 85428 58492
rect 85260 57598 85262 57650
rect 85314 57598 85316 57650
rect 85260 57586 85316 57598
rect 85148 56642 85204 56654
rect 85148 56590 85150 56642
rect 85202 56590 85204 56642
rect 85148 55300 85204 56590
rect 85484 56308 85540 60956
rect 85820 60946 85876 60958
rect 85596 60786 85652 60798
rect 85596 60734 85598 60786
rect 85650 60734 85652 60786
rect 85596 60564 85652 60734
rect 85596 60498 85652 60508
rect 85708 60788 85764 60798
rect 85596 60004 85652 60014
rect 85596 59910 85652 59948
rect 85708 59108 85764 60732
rect 86044 60004 86100 60014
rect 86044 59910 86100 59948
rect 86156 59892 86212 61516
rect 86604 61516 86772 61572
rect 86828 62580 86884 62590
rect 86380 60786 86436 60798
rect 86380 60734 86382 60786
rect 86434 60734 86436 60786
rect 86268 59892 86324 59902
rect 86156 59890 86324 59892
rect 86156 59838 86270 59890
rect 86322 59838 86324 59890
rect 86156 59836 86324 59838
rect 86268 59826 86324 59836
rect 86380 59892 86436 60734
rect 86604 60676 86660 61516
rect 86716 61348 86772 61358
rect 86828 61348 86884 62524
rect 86716 61346 86884 61348
rect 86716 61294 86718 61346
rect 86770 61294 86884 61346
rect 86716 61292 86884 61294
rect 86716 61282 86772 61292
rect 87052 61124 87108 63644
rect 87388 63140 87444 63868
rect 87388 63084 87556 63140
rect 87388 62916 87444 62926
rect 87276 62914 87444 62916
rect 87276 62862 87390 62914
rect 87442 62862 87444 62914
rect 87276 62860 87444 62862
rect 87276 62692 87332 62860
rect 87388 62850 87444 62860
rect 87276 62466 87332 62636
rect 87276 62414 87278 62466
rect 87330 62414 87332 62466
rect 87276 62402 87332 62414
rect 87500 62466 87556 63084
rect 87612 62578 87668 63980
rect 87724 63812 87780 65324
rect 87948 64706 88004 66220
rect 88060 65716 88116 65726
rect 88060 65622 88116 65660
rect 88284 65604 88340 66894
rect 88844 66164 88900 68348
rect 88284 65538 88340 65548
rect 88620 66108 88900 66164
rect 88956 67956 89012 67966
rect 88172 65492 88228 65502
rect 88172 65398 88228 65436
rect 88620 65380 88676 66108
rect 88844 65828 88900 65838
rect 88620 65324 88788 65380
rect 88060 65268 88116 65278
rect 88060 65266 88676 65268
rect 88060 65214 88062 65266
rect 88114 65214 88676 65266
rect 88060 65212 88676 65214
rect 88060 65202 88116 65212
rect 87948 64654 87950 64706
rect 88002 64654 88004 64706
rect 87948 64642 88004 64654
rect 88508 65044 88564 65054
rect 88396 64596 88452 64606
rect 88396 64146 88452 64540
rect 88396 64094 88398 64146
rect 88450 64094 88452 64146
rect 87948 63812 88004 63822
rect 87724 63810 88004 63812
rect 87724 63758 87950 63810
rect 88002 63758 88004 63810
rect 87724 63756 88004 63758
rect 87948 62692 88004 63756
rect 88396 63364 88452 64094
rect 88396 63298 88452 63308
rect 88396 63140 88452 63150
rect 88284 63084 88396 63140
rect 87948 62626 88004 62636
rect 88060 63026 88116 63038
rect 88060 62974 88062 63026
rect 88114 62974 88116 63026
rect 88060 62916 88116 62974
rect 87612 62526 87614 62578
rect 87666 62526 87668 62578
rect 87612 62514 87668 62526
rect 87500 62414 87502 62466
rect 87554 62414 87556 62466
rect 87500 62402 87556 62414
rect 87836 62468 87892 62478
rect 87836 62374 87892 62412
rect 87612 61684 87668 61694
rect 87612 61590 87668 61628
rect 87164 61348 87220 61358
rect 87164 61254 87220 61292
rect 87052 61068 87220 61124
rect 87052 60788 87108 60798
rect 87052 60694 87108 60732
rect 86604 60610 86660 60620
rect 86716 59892 86772 59902
rect 86380 59890 86772 59892
rect 86380 59838 86718 59890
rect 86770 59838 86772 59890
rect 86380 59836 86772 59838
rect 86380 59108 86436 59836
rect 86716 59826 86772 59836
rect 85708 59106 85876 59108
rect 85708 59054 85710 59106
rect 85762 59054 85876 59106
rect 85708 59052 85876 59054
rect 85708 59042 85764 59052
rect 85372 56252 85540 56308
rect 85260 55300 85316 55310
rect 85204 55298 85316 55300
rect 85204 55246 85262 55298
rect 85314 55246 85316 55298
rect 85204 55244 85316 55246
rect 85148 55234 85204 55244
rect 85260 55234 85316 55244
rect 85260 54628 85316 54638
rect 85260 54534 85316 54572
rect 84700 54404 84756 54414
rect 84700 54310 84756 54348
rect 85148 53620 85204 53630
rect 85148 53526 85204 53564
rect 85260 52836 85316 52846
rect 85260 52742 85316 52780
rect 84924 51268 84980 51278
rect 84588 50082 84644 50092
rect 84812 50596 84868 50606
rect 84812 50036 84868 50540
rect 84812 49970 84868 49980
rect 84140 47518 84142 47570
rect 84194 47518 84196 47570
rect 84140 47506 84196 47518
rect 84364 48524 84532 48580
rect 84588 48916 84644 48926
rect 83132 46900 83188 46910
rect 83132 46004 83188 46844
rect 83916 46004 83972 46014
rect 83132 46002 83972 46004
rect 83132 45950 83918 46002
rect 83970 45950 83972 46002
rect 83132 45948 83972 45950
rect 83132 45778 83188 45948
rect 83916 45938 83972 45948
rect 83132 45726 83134 45778
rect 83186 45726 83188 45778
rect 83132 45714 83188 45726
rect 84252 45892 84308 45902
rect 83356 45668 83412 45678
rect 83244 41076 83300 41086
rect 83244 40982 83300 41020
rect 82908 39666 82964 39676
rect 82348 39526 82404 39564
rect 82460 39564 82740 39620
rect 83244 39620 83300 39630
rect 82460 38836 82516 39564
rect 83244 39526 83300 39564
rect 82572 39396 82628 39406
rect 82572 39394 83300 39396
rect 82572 39342 82574 39394
rect 82626 39342 83300 39394
rect 82572 39340 83300 39342
rect 82572 39330 82628 39340
rect 82124 37940 82180 37950
rect 81900 37938 82180 37940
rect 81900 37886 82126 37938
rect 82178 37886 82180 37938
rect 81900 37884 82180 37886
rect 81900 37490 81956 37884
rect 82124 37874 82180 37884
rect 81900 37438 81902 37490
rect 81954 37438 81956 37490
rect 81900 37426 81956 37438
rect 82236 37268 82292 37278
rect 82236 37174 82292 37212
rect 81788 35924 81844 36764
rect 82460 36596 82516 38780
rect 82572 39060 82628 39070
rect 82572 38834 82628 39004
rect 83244 38946 83300 39340
rect 83244 38894 83246 38946
rect 83298 38894 83300 38946
rect 83244 38882 83300 38894
rect 82572 38782 82574 38834
rect 82626 38782 82628 38834
rect 82572 38770 82628 38782
rect 83244 38164 83300 38174
rect 82908 37268 82964 37278
rect 82908 37174 82964 37212
rect 83244 37266 83300 38108
rect 83244 37214 83246 37266
rect 83298 37214 83300 37266
rect 83244 37202 83300 37214
rect 83356 36708 83412 45612
rect 84252 44994 84308 45836
rect 84252 44942 84254 44994
rect 84306 44942 84308 44994
rect 84252 44930 84308 44942
rect 83916 44322 83972 44334
rect 83916 44270 83918 44322
rect 83970 44270 83972 44322
rect 83916 42084 83972 44270
rect 83804 40962 83860 40974
rect 83804 40910 83806 40962
rect 83858 40910 83860 40962
rect 83804 40292 83860 40910
rect 83916 40404 83972 42028
rect 83916 40272 83972 40348
rect 84140 42644 84196 42654
rect 83804 39732 83860 40236
rect 83804 39666 83860 39676
rect 84140 40180 84196 42588
rect 84252 41860 84308 41870
rect 84364 41860 84420 48524
rect 84476 48132 84532 48142
rect 84588 48132 84644 48860
rect 84476 48130 84644 48132
rect 84476 48078 84478 48130
rect 84530 48078 84644 48130
rect 84476 48076 84644 48078
rect 84476 48066 84532 48076
rect 84476 47572 84532 47582
rect 84476 47478 84532 47516
rect 84476 45780 84532 45790
rect 84476 45686 84532 45724
rect 84924 45668 84980 51212
rect 85260 50484 85316 50522
rect 85260 50418 85316 50428
rect 85036 50036 85092 50046
rect 85372 50036 85428 56252
rect 85596 55188 85652 55198
rect 85596 54738 85652 55132
rect 85596 54686 85598 54738
rect 85650 54686 85652 54738
rect 85596 54674 85652 54686
rect 85484 52164 85540 52174
rect 85484 50428 85540 52108
rect 85708 51940 85764 51950
rect 85708 51266 85764 51884
rect 85708 51214 85710 51266
rect 85762 51214 85764 51266
rect 85484 50372 85652 50428
rect 85036 50034 85428 50036
rect 85036 49982 85038 50034
rect 85090 49982 85428 50034
rect 85036 49980 85428 49982
rect 85036 49812 85092 49980
rect 85036 49746 85092 49756
rect 85260 49700 85316 49710
rect 85484 49700 85540 49710
rect 85316 49698 85540 49700
rect 85316 49646 85486 49698
rect 85538 49646 85540 49698
rect 85316 49644 85540 49646
rect 85036 48916 85092 48926
rect 85036 48130 85092 48860
rect 85036 48078 85038 48130
rect 85090 48078 85092 48130
rect 85036 48066 85092 48078
rect 85148 47684 85204 47694
rect 85148 46898 85204 47628
rect 85148 46846 85150 46898
rect 85202 46846 85204 46898
rect 85148 46834 85204 46846
rect 84924 45602 84980 45612
rect 84924 45106 84980 45118
rect 84924 45054 84926 45106
rect 84978 45054 84980 45106
rect 84700 43426 84756 43438
rect 84700 43374 84702 43426
rect 84754 43374 84756 43426
rect 84700 42084 84756 43374
rect 84700 42018 84756 42028
rect 84252 41858 84420 41860
rect 84252 41806 84254 41858
rect 84306 41806 84420 41858
rect 84252 41804 84420 41806
rect 84924 41970 84980 45054
rect 85260 43708 85316 49644
rect 85484 49634 85540 49644
rect 85596 49700 85652 50372
rect 85596 49634 85652 49644
rect 85708 49252 85764 51214
rect 85820 50708 85876 59052
rect 86380 59042 86436 59052
rect 86492 58212 86548 58222
rect 85932 57652 85988 57662
rect 85932 57558 85988 57596
rect 85932 55300 85988 55310
rect 85932 54740 85988 55244
rect 86044 55188 86100 55198
rect 86044 55094 86100 55132
rect 86044 54740 86100 54750
rect 85932 54738 86100 54740
rect 85932 54686 86046 54738
rect 86098 54686 86100 54738
rect 85932 54684 86100 54686
rect 86044 54674 86100 54684
rect 86380 53620 86436 53630
rect 86380 53526 86436 53564
rect 86044 53508 86100 53518
rect 86044 52836 86100 53452
rect 86044 52274 86100 52780
rect 86044 52222 86046 52274
rect 86098 52222 86100 52274
rect 86044 52210 86100 52222
rect 86380 52162 86436 52174
rect 86380 52110 86382 52162
rect 86434 52110 86436 52162
rect 86380 51940 86436 52110
rect 86380 51874 86436 51884
rect 85820 50652 85988 50708
rect 85820 50482 85876 50494
rect 85820 50430 85822 50482
rect 85874 50430 85876 50482
rect 85820 50372 85876 50430
rect 85820 49476 85876 50316
rect 85820 49410 85876 49420
rect 85932 49252 85988 50652
rect 86492 50260 86548 58156
rect 86828 58212 86884 58222
rect 86828 58210 86996 58212
rect 86828 58158 86830 58210
rect 86882 58158 86996 58210
rect 86828 58156 86996 58158
rect 86828 58146 86884 58156
rect 86828 57650 86884 57662
rect 86828 57598 86830 57650
rect 86882 57598 86884 57650
rect 86828 57428 86884 57598
rect 86828 57362 86884 57372
rect 86940 57316 86996 58156
rect 86268 50204 86548 50260
rect 86604 56308 86660 56318
rect 85708 49196 85876 49252
rect 85932 49196 86100 49252
rect 85596 49028 85652 49066
rect 85596 48962 85652 48972
rect 85708 48916 85764 48926
rect 85708 48822 85764 48860
rect 85820 47684 85876 49196
rect 85932 49028 85988 49038
rect 85932 48934 85988 48972
rect 85820 47618 85876 47628
rect 85484 47460 85540 47470
rect 85484 46564 85540 47404
rect 85596 47458 85652 47470
rect 85596 47406 85598 47458
rect 85650 47406 85652 47458
rect 85596 46788 85652 47406
rect 86044 47236 86100 49196
rect 86268 49138 86324 50204
rect 86492 49924 86548 49934
rect 86492 49830 86548 49868
rect 86268 49086 86270 49138
rect 86322 49086 86324 49138
rect 86268 48916 86324 49086
rect 86380 49810 86436 49822
rect 86380 49758 86382 49810
rect 86434 49758 86436 49810
rect 86380 49028 86436 49758
rect 86380 48962 86436 48972
rect 86268 48850 86324 48860
rect 86492 48132 86548 48142
rect 86492 47458 86548 48076
rect 86492 47406 86494 47458
rect 86546 47406 86548 47458
rect 86492 47394 86548 47406
rect 86044 47170 86100 47180
rect 85596 46722 85652 46732
rect 86268 46788 86324 46798
rect 85596 46564 85652 46574
rect 85484 46562 85652 46564
rect 85484 46510 85598 46562
rect 85650 46510 85652 46562
rect 85484 46508 85652 46510
rect 85596 46498 85652 46508
rect 85708 45892 85764 45902
rect 85708 45798 85764 45836
rect 85932 45780 85988 45790
rect 85932 45686 85988 45724
rect 86268 45780 86324 46732
rect 85372 45666 85428 45678
rect 85372 45614 85374 45666
rect 85426 45614 85428 45666
rect 86268 45648 86324 45724
rect 85372 44322 85428 45614
rect 85372 44270 85374 44322
rect 85426 44270 85428 44322
rect 85372 44258 85428 44270
rect 85596 44994 85652 45006
rect 85596 44942 85598 44994
rect 85650 44942 85652 44994
rect 85596 44210 85652 44942
rect 85596 44158 85598 44210
rect 85650 44158 85652 44210
rect 85596 44146 85652 44158
rect 84924 41918 84926 41970
rect 84978 41918 84980 41970
rect 84252 41298 84308 41804
rect 84252 41246 84254 41298
rect 84306 41246 84308 41298
rect 84252 41076 84308 41246
rect 84252 41010 84308 41020
rect 84924 40292 84980 41918
rect 84924 40226 84980 40236
rect 85148 43652 85316 43708
rect 83580 39618 83636 39630
rect 84140 39620 84196 40124
rect 85148 39732 85204 43652
rect 86156 42756 86212 42766
rect 86156 42662 86212 42700
rect 85260 42644 85316 42654
rect 85260 42550 85316 42588
rect 86380 42644 86436 42654
rect 86380 42550 86436 42588
rect 85820 42530 85876 42542
rect 85820 42478 85822 42530
rect 85874 42478 85876 42530
rect 85596 41858 85652 41870
rect 85596 41806 85598 41858
rect 85650 41806 85652 41858
rect 85596 41074 85652 41806
rect 85820 41186 85876 42478
rect 86604 42532 86660 56252
rect 86828 54516 86884 54526
rect 86828 54422 86884 54460
rect 86940 53620 86996 57260
rect 86940 53526 86996 53564
rect 87052 53508 87108 53518
rect 87052 53414 87108 53452
rect 86940 52162 86996 52174
rect 86940 52110 86942 52162
rect 86994 52110 86996 52162
rect 86940 51940 86996 52110
rect 87052 52052 87108 52062
rect 87164 52052 87220 61068
rect 87948 60786 88004 60798
rect 87948 60734 87950 60786
rect 88002 60734 88004 60786
rect 87948 60564 88004 60734
rect 87948 60498 88004 60508
rect 88060 60340 88116 62860
rect 87948 60284 88116 60340
rect 88172 62692 88228 62702
rect 87500 60002 87556 60014
rect 87500 59950 87502 60002
rect 87554 59950 87556 60002
rect 87500 59444 87556 59950
rect 87500 59378 87556 59388
rect 87724 58322 87780 58334
rect 87724 58270 87726 58322
rect 87778 58270 87780 58322
rect 87276 58212 87332 58222
rect 87276 58118 87332 58156
rect 87500 57652 87556 57662
rect 87500 57540 87556 57596
rect 87500 57538 87668 57540
rect 87500 57486 87502 57538
rect 87554 57486 87668 57538
rect 87500 57484 87668 57486
rect 87500 57474 87556 57484
rect 87388 57204 87444 57214
rect 87388 56978 87444 57148
rect 87388 56926 87390 56978
rect 87442 56926 87444 56978
rect 87388 56914 87444 56926
rect 87500 56084 87556 56094
rect 87500 55990 87556 56028
rect 87500 54740 87556 54750
rect 87500 54646 87556 54684
rect 87388 54516 87444 54526
rect 87276 54514 87444 54516
rect 87276 54462 87390 54514
rect 87442 54462 87444 54514
rect 87276 54460 87444 54462
rect 87276 53730 87332 54460
rect 87388 54450 87444 54460
rect 87276 53678 87278 53730
rect 87330 53678 87332 53730
rect 87276 53666 87332 53678
rect 87500 54290 87556 54302
rect 87500 54238 87502 54290
rect 87554 54238 87556 54290
rect 87388 53060 87444 53070
rect 87500 53060 87556 54238
rect 87388 53058 87556 53060
rect 87388 53006 87390 53058
rect 87442 53006 87556 53058
rect 87388 53004 87556 53006
rect 87388 52994 87444 53004
rect 87500 52164 87556 52174
rect 87500 52070 87556 52108
rect 87052 52050 87220 52052
rect 87052 51998 87054 52050
rect 87106 51998 87220 52050
rect 87052 51996 87220 51998
rect 87052 51986 87108 51996
rect 86940 51874 86996 51884
rect 87276 50482 87332 50494
rect 87276 50430 87278 50482
rect 87330 50430 87332 50482
rect 87276 50372 87332 50430
rect 86716 49812 86772 49822
rect 87276 49812 87332 50316
rect 87612 50148 87668 57484
rect 87724 57316 87780 58270
rect 87836 58324 87892 58334
rect 87836 58230 87892 58268
rect 87948 58100 88004 60284
rect 88172 59332 88228 62636
rect 88284 62242 88340 63084
rect 88396 63008 88452 63084
rect 88284 62190 88286 62242
rect 88338 62190 88340 62242
rect 88284 61572 88340 62190
rect 88284 61506 88340 61516
rect 88508 61010 88564 64988
rect 88620 64818 88676 65212
rect 88620 64766 88622 64818
rect 88674 64766 88676 64818
rect 88620 64754 88676 64766
rect 88620 64372 88676 64382
rect 88620 62356 88676 64316
rect 88732 63252 88788 65324
rect 88732 63186 88788 63196
rect 88844 63138 88900 65772
rect 88956 65604 89012 67900
rect 89516 67228 89572 68684
rect 89628 68738 89684 69916
rect 89628 68686 89630 68738
rect 89682 68686 89684 68738
rect 89628 68674 89684 68686
rect 89068 67172 89124 67182
rect 89068 65828 89124 67116
rect 89068 65762 89124 65772
rect 89292 67172 89572 67228
rect 88956 65538 89012 65548
rect 89180 65492 89236 65502
rect 89180 65398 89236 65436
rect 89292 64148 89348 67172
rect 89404 65602 89460 65614
rect 89404 65550 89406 65602
rect 89458 65550 89460 65602
rect 89404 64820 89460 65550
rect 89516 65604 89572 65614
rect 89516 65510 89572 65548
rect 89404 64754 89460 64764
rect 89180 64092 89348 64148
rect 88844 63086 88846 63138
rect 88898 63086 88900 63138
rect 88844 63074 88900 63086
rect 88956 63364 89012 63374
rect 88620 62290 88676 62300
rect 88844 61684 88900 61694
rect 88956 61684 89012 63308
rect 89068 62914 89124 62926
rect 89068 62862 89070 62914
rect 89122 62862 89124 62914
rect 89068 62468 89124 62862
rect 89068 62402 89124 62412
rect 89180 62244 89236 64092
rect 89292 63924 89348 63934
rect 89292 63830 89348 63868
rect 89628 63922 89684 63934
rect 89628 63870 89630 63922
rect 89682 63870 89684 63922
rect 89516 63700 89572 63710
rect 89516 63364 89572 63644
rect 89516 63138 89572 63308
rect 89516 63086 89518 63138
rect 89570 63086 89572 63138
rect 89516 63074 89572 63086
rect 89628 63140 89684 63870
rect 89628 63074 89684 63084
rect 89292 62468 89348 62478
rect 89292 62374 89348 62412
rect 88844 61682 89012 61684
rect 88844 61630 88846 61682
rect 88898 61630 89012 61682
rect 88844 61628 89012 61630
rect 89068 62188 89236 62244
rect 89516 62356 89572 62366
rect 89628 62356 89684 62366
rect 89572 62354 89684 62356
rect 89572 62302 89630 62354
rect 89682 62302 89684 62354
rect 89572 62300 89684 62302
rect 88844 61618 88900 61628
rect 88508 60958 88510 61010
rect 88562 60958 88564 61010
rect 88508 60676 88564 60958
rect 88508 60610 88564 60620
rect 89068 60114 89124 62188
rect 89180 61684 89236 61694
rect 89516 61684 89572 62300
rect 89628 62290 89684 62300
rect 89180 61682 89572 61684
rect 89180 61630 89182 61682
rect 89234 61630 89572 61682
rect 89180 61628 89572 61630
rect 89180 61618 89236 61628
rect 89628 61572 89684 61582
rect 89628 61478 89684 61516
rect 89740 61348 89796 70140
rect 89852 63140 89908 70924
rect 90860 70914 90916 70924
rect 91308 71092 91364 71102
rect 91308 70978 91364 71036
rect 91308 70926 91310 70978
rect 91362 70926 91364 70978
rect 91308 70914 91364 70926
rect 91196 70868 91252 70878
rect 90972 70866 91252 70868
rect 90972 70814 91198 70866
rect 91250 70814 91252 70866
rect 90972 70812 91252 70814
rect 90300 70306 90356 70318
rect 90300 70254 90302 70306
rect 90354 70254 90356 70306
rect 90188 70196 90244 70206
rect 89964 70194 90244 70196
rect 89964 70142 90190 70194
rect 90242 70142 90244 70194
rect 89964 70140 90244 70142
rect 89964 65490 90020 70140
rect 90188 70130 90244 70140
rect 90300 69412 90356 70254
rect 90524 70196 90580 70206
rect 90524 70194 90692 70196
rect 90524 70142 90526 70194
rect 90578 70142 90692 70194
rect 90524 70140 90692 70142
rect 90524 70130 90580 70140
rect 90300 69346 90356 69356
rect 90524 68964 90580 68974
rect 90524 68850 90580 68908
rect 90524 68798 90526 68850
rect 90578 68798 90580 68850
rect 90524 68786 90580 68798
rect 90188 68740 90244 68750
rect 90188 68626 90244 68684
rect 90188 68574 90190 68626
rect 90242 68574 90244 68626
rect 90188 68404 90244 68574
rect 90188 68338 90244 68348
rect 90636 67956 90692 70140
rect 90972 70082 91028 70812
rect 91196 70802 91252 70812
rect 90972 70030 90974 70082
rect 91026 70030 91028 70082
rect 90972 69972 91028 70030
rect 90972 69906 91028 69916
rect 91196 68628 91252 68638
rect 91196 68534 91252 68572
rect 90972 68068 91028 68078
rect 90860 67956 90916 67966
rect 90636 67954 90916 67956
rect 90636 67902 90862 67954
rect 90914 67902 90916 67954
rect 90636 67900 90916 67902
rect 90860 67890 90916 67900
rect 90860 67060 90916 67070
rect 90860 66498 90916 67004
rect 90860 66446 90862 66498
rect 90914 66446 90916 66498
rect 90860 66434 90916 66446
rect 90188 66388 90244 66398
rect 89964 65438 89966 65490
rect 90018 65438 90020 65490
rect 89964 65426 90020 65438
rect 90076 66386 90244 66388
rect 90076 66334 90190 66386
rect 90242 66334 90244 66386
rect 90076 66332 90244 66334
rect 90076 66052 90132 66332
rect 90188 66322 90244 66332
rect 90972 66388 91028 68012
rect 91420 67228 91476 74284
rect 91644 74228 91700 74238
rect 91644 74134 91700 74172
rect 91756 73332 91812 73342
rect 91756 73238 91812 73276
rect 91756 72436 91812 72446
rect 91644 69300 91700 69310
rect 91644 69206 91700 69244
rect 90972 66322 91028 66332
rect 91196 67172 91476 67228
rect 91532 67842 91588 67854
rect 91532 67790 91534 67842
rect 91586 67790 91588 67842
rect 90972 66164 91028 66174
rect 90076 63922 90132 65996
rect 90860 66052 90916 66062
rect 90860 65958 90916 65996
rect 90188 65828 90244 65838
rect 90188 65714 90244 65772
rect 90188 65662 90190 65714
rect 90242 65662 90244 65714
rect 90188 65650 90244 65662
rect 90860 65716 90916 65726
rect 90972 65716 91028 66108
rect 90916 65660 91028 65716
rect 90300 65604 90356 65614
rect 90300 65510 90356 65548
rect 90636 65604 90692 65614
rect 90860 65584 90916 65660
rect 90076 63870 90078 63922
rect 90130 63870 90132 63922
rect 90076 63858 90132 63870
rect 90188 64820 90244 64830
rect 90076 63252 90132 63262
rect 90076 63140 90132 63196
rect 89852 63138 90132 63140
rect 89852 63086 90078 63138
rect 90130 63086 90132 63138
rect 89852 63084 90132 63086
rect 90076 63074 90132 63084
rect 90188 62354 90244 64764
rect 90300 64148 90356 64158
rect 90300 64054 90356 64092
rect 90412 63924 90468 63934
rect 90300 63028 90356 63038
rect 90300 62578 90356 62972
rect 90300 62526 90302 62578
rect 90354 62526 90356 62578
rect 90300 62514 90356 62526
rect 90188 62302 90190 62354
rect 90242 62302 90244 62354
rect 90188 62290 90244 62302
rect 89740 61292 89908 61348
rect 89740 60788 89796 60798
rect 89740 60694 89796 60732
rect 89292 60674 89348 60686
rect 89292 60622 89294 60674
rect 89346 60622 89348 60674
rect 89292 60564 89348 60622
rect 89852 60564 89908 61292
rect 89292 60498 89348 60508
rect 89740 60508 89908 60564
rect 89068 60062 89070 60114
rect 89122 60062 89124 60114
rect 88396 60002 88452 60014
rect 88396 59950 88398 60002
rect 88450 59950 88452 60002
rect 88396 59780 88452 59950
rect 89068 60004 89124 60062
rect 89068 59938 89124 59948
rect 88396 59714 88452 59724
rect 88844 59780 88900 59790
rect 88172 59266 88228 59276
rect 88508 58548 88564 58558
rect 88564 58492 88788 58548
rect 88508 58454 88564 58492
rect 88060 58212 88116 58222
rect 88060 58210 88340 58212
rect 88060 58158 88062 58210
rect 88114 58158 88340 58210
rect 88060 58156 88340 58158
rect 88060 58146 88116 58156
rect 87724 57250 87780 57260
rect 87836 58044 88004 58100
rect 87836 55468 87892 58044
rect 88284 57762 88340 58156
rect 88284 57710 88286 57762
rect 88338 57710 88340 57762
rect 88284 57698 88340 57710
rect 88396 57762 88452 57774
rect 88396 57710 88398 57762
rect 88450 57710 88452 57762
rect 88172 57428 88228 57438
rect 87948 57316 88004 57326
rect 87948 56978 88004 57260
rect 87948 56926 87950 56978
rect 88002 56926 88004 56978
rect 87948 56914 88004 56926
rect 86716 49810 87220 49812
rect 86716 49758 86718 49810
rect 86770 49758 87220 49810
rect 86716 49756 87220 49758
rect 86716 49746 86772 49756
rect 86940 49588 86996 49598
rect 86940 47458 86996 49532
rect 87164 48354 87220 49756
rect 87276 49746 87332 49756
rect 87388 50092 87668 50148
rect 87724 55412 87892 55468
rect 87164 48302 87166 48354
rect 87218 48302 87220 48354
rect 87164 48290 87220 48302
rect 86940 47406 86942 47458
rect 86994 47406 86996 47458
rect 86940 47394 86996 47406
rect 87388 42868 87444 50092
rect 87612 49922 87668 49934
rect 87612 49870 87614 49922
rect 87666 49870 87668 49922
rect 87500 49812 87556 49822
rect 87500 49718 87556 49756
rect 87612 47460 87668 49870
rect 87724 48020 87780 55412
rect 88172 55410 88228 57372
rect 88396 56532 88452 57710
rect 88620 57652 88676 57662
rect 88620 57558 88676 57596
rect 88508 57316 88564 57326
rect 88508 56866 88564 57260
rect 88620 57204 88676 57214
rect 88620 57090 88676 57148
rect 88620 57038 88622 57090
rect 88674 57038 88676 57090
rect 88620 57026 88676 57038
rect 88508 56814 88510 56866
rect 88562 56814 88564 56866
rect 88508 56802 88564 56814
rect 88620 56756 88676 56766
rect 88732 56756 88788 58492
rect 88620 56754 88788 56756
rect 88620 56702 88622 56754
rect 88674 56702 88788 56754
rect 88620 56700 88788 56702
rect 88620 56690 88676 56700
rect 88284 56476 88452 56532
rect 88284 56196 88340 56476
rect 88620 56308 88676 56318
rect 88620 56214 88676 56252
rect 88284 56102 88340 56140
rect 88396 56196 88452 56206
rect 88396 56194 88564 56196
rect 88396 56142 88398 56194
rect 88450 56142 88564 56194
rect 88396 56140 88564 56142
rect 88396 56130 88452 56140
rect 88172 55358 88174 55410
rect 88226 55358 88228 55410
rect 88172 55346 88228 55358
rect 88508 54738 88564 56140
rect 88508 54686 88510 54738
rect 88562 54686 88564 54738
rect 88508 54674 88564 54686
rect 87836 54628 87892 54638
rect 87836 53842 87892 54572
rect 88284 54626 88340 54638
rect 88284 54574 88286 54626
rect 88338 54574 88340 54626
rect 88172 54516 88228 54526
rect 88172 54422 88228 54460
rect 88284 54292 88340 54574
rect 88284 54226 88340 54236
rect 87836 53790 87838 53842
rect 87890 53790 87892 53842
rect 87836 53778 87892 53790
rect 88172 52946 88228 52958
rect 88172 52894 88174 52946
rect 88226 52894 88228 52946
rect 87836 49812 87892 49822
rect 87836 49718 87892 49756
rect 87724 47954 87780 47964
rect 87836 49588 87892 49598
rect 87724 47460 87780 47470
rect 87612 47404 87724 47460
rect 87724 47366 87780 47404
rect 87612 47236 87668 47246
rect 87612 47142 87668 47180
rect 87724 46788 87780 46798
rect 87836 46788 87892 49532
rect 88172 49140 88228 52894
rect 88284 52162 88340 52174
rect 88284 52110 88286 52162
rect 88338 52110 88340 52162
rect 88284 50036 88340 52110
rect 88284 49970 88340 49980
rect 88396 49924 88452 49934
rect 88396 49922 88564 49924
rect 88396 49870 88398 49922
rect 88450 49870 88564 49922
rect 88396 49868 88564 49870
rect 88396 49858 88452 49868
rect 88284 49812 88340 49822
rect 88284 49718 88340 49756
rect 88396 49588 88452 49598
rect 88396 49494 88452 49532
rect 87948 49138 88228 49140
rect 87948 49086 88174 49138
rect 88226 49086 88228 49138
rect 87948 49084 88228 49086
rect 87948 48244 88004 49084
rect 88172 49074 88228 49084
rect 87948 48242 88452 48244
rect 87948 48190 87950 48242
rect 88002 48190 88452 48242
rect 87948 48188 88452 48190
rect 87948 48178 88004 48188
rect 87724 46786 87892 46788
rect 87724 46734 87726 46786
rect 87778 46734 87892 46786
rect 87724 46732 87892 46734
rect 88060 48020 88116 48030
rect 87724 46722 87780 46732
rect 87724 45780 87780 45790
rect 87724 44994 87780 45724
rect 87724 44942 87726 44994
rect 87778 44942 87780 44994
rect 87724 44930 87780 44942
rect 87500 42868 87556 42878
rect 86940 42866 87780 42868
rect 86940 42814 87502 42866
rect 87554 42814 87780 42866
rect 86940 42812 87780 42814
rect 86604 42466 86660 42476
rect 86716 42756 86772 42766
rect 86716 41298 86772 42700
rect 86940 42642 86996 42812
rect 87500 42802 87556 42812
rect 86940 42590 86942 42642
rect 86994 42590 86996 42642
rect 86940 42578 86996 42590
rect 87724 41858 87780 42812
rect 87724 41806 87726 41858
rect 87778 41806 87780 41858
rect 87724 41794 87780 41806
rect 86716 41246 86718 41298
rect 86770 41246 86772 41298
rect 86716 41234 86772 41246
rect 85820 41134 85822 41186
rect 85874 41134 85876 41186
rect 85820 41122 85876 41134
rect 85596 41022 85598 41074
rect 85650 41022 85652 41074
rect 85596 41010 85652 41022
rect 85820 40292 85876 40302
rect 83580 39566 83582 39618
rect 83634 39566 83636 39618
rect 83580 38164 83636 39566
rect 83580 38098 83636 38108
rect 83916 39618 84196 39620
rect 83916 39566 84142 39618
rect 84194 39566 84196 39618
rect 83916 39564 84196 39566
rect 83132 36652 83412 36708
rect 83804 37378 83860 37390
rect 83804 37326 83806 37378
rect 83858 37326 83860 37378
rect 83804 37156 83860 37326
rect 83916 37266 83972 39564
rect 84140 39554 84196 39564
rect 84364 39730 85428 39732
rect 84364 39678 85150 39730
rect 85202 39678 85428 39730
rect 84364 39676 85428 39678
rect 84364 39506 84420 39676
rect 85148 39666 85204 39676
rect 84364 39454 84366 39506
rect 84418 39454 84420 39506
rect 84364 39442 84420 39454
rect 84476 39060 84532 39070
rect 84252 38164 84308 38174
rect 84252 38070 84308 38108
rect 83916 37214 83918 37266
rect 83970 37214 83972 37266
rect 83916 37202 83972 37214
rect 82572 36596 82628 36606
rect 82460 36594 82628 36596
rect 82460 36542 82574 36594
rect 82626 36542 82628 36594
rect 82460 36540 82628 36542
rect 82572 36530 82628 36540
rect 81788 35364 81844 35868
rect 82460 35924 82516 35934
rect 83132 35924 83188 36652
rect 82460 35922 83188 35924
rect 82460 35870 82462 35922
rect 82514 35870 83188 35922
rect 82460 35868 83188 35870
rect 82460 35858 82516 35868
rect 81788 35298 81844 35308
rect 81676 34974 81678 35026
rect 81730 34974 81732 35026
rect 81676 34804 81732 34974
rect 81676 34738 81732 34748
rect 82124 34916 82180 34926
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 81116 33684 81172 33694
rect 81116 33458 81172 33628
rect 82124 33684 82180 34860
rect 82348 34690 82404 34702
rect 82348 34638 82350 34690
rect 82402 34638 82404 34690
rect 82348 34244 82404 34638
rect 82348 34178 82404 34188
rect 82124 33570 82180 33628
rect 82124 33518 82126 33570
rect 82178 33518 82180 33570
rect 82124 33506 82180 33518
rect 82460 34132 82516 34142
rect 82460 34018 82516 34076
rect 82460 33966 82462 34018
rect 82514 33966 82516 34018
rect 81116 33406 81118 33458
rect 81170 33406 81172 33458
rect 81116 33394 81172 33406
rect 81788 33122 81844 33134
rect 81788 33070 81790 33122
rect 81842 33070 81844 33122
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 81340 32788 81396 32798
rect 81340 32694 81396 32732
rect 81676 32676 81732 32686
rect 81788 32676 81844 33070
rect 81676 32674 81844 32676
rect 81676 32622 81678 32674
rect 81730 32622 81844 32674
rect 81676 32620 81844 32622
rect 81676 32610 81732 32620
rect 82348 32564 82404 32574
rect 82460 32564 82516 33966
rect 82348 32562 82516 32564
rect 82348 32510 82350 32562
rect 82402 32510 82516 32562
rect 82348 32508 82516 32510
rect 77420 31892 77588 31948
rect 81004 31892 81956 31948
rect 76972 25218 77028 25228
rect 73388 12674 73444 12684
rect 69132 3332 69188 3342
rect 69132 3238 69188 3276
rect 77532 2884 77588 31892
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 81276 25116 81540 25126
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 81900 8428 81956 31892
rect 82348 30996 82404 32508
rect 82348 30930 82404 30940
rect 82572 8428 82628 35868
rect 83132 35698 83188 35868
rect 83132 35646 83134 35698
rect 83186 35646 83188 35698
rect 83132 35634 83188 35646
rect 83356 35812 83412 35822
rect 83804 35812 83860 37100
rect 83356 35810 83860 35812
rect 83356 35758 83358 35810
rect 83410 35758 83860 35810
rect 83356 35756 83860 35758
rect 84476 35922 84532 39004
rect 85148 39060 85204 39070
rect 85148 38162 85204 39004
rect 85372 38722 85428 39676
rect 85820 39060 85876 40236
rect 87948 39732 88004 39742
rect 87948 39638 88004 39676
rect 85820 38928 85876 39004
rect 85372 38670 85374 38722
rect 85426 38670 85428 38722
rect 85372 38658 85428 38670
rect 85148 38110 85150 38162
rect 85202 38110 85204 38162
rect 85148 38098 85204 38110
rect 84588 37156 84644 37166
rect 84588 37062 84644 37100
rect 86716 36596 86772 36606
rect 84476 35870 84478 35922
rect 84530 35870 84532 35922
rect 82908 35252 82964 35262
rect 82684 34916 82740 34926
rect 82684 34822 82740 34860
rect 82908 34804 82964 35196
rect 82796 34802 82964 34804
rect 82796 34750 82910 34802
rect 82962 34750 82964 34802
rect 82796 34748 82964 34750
rect 82796 33348 82852 34748
rect 82908 34738 82964 34748
rect 83244 34804 83300 34814
rect 83244 34710 83300 34748
rect 82796 33216 82852 33292
rect 82908 33236 82964 33246
rect 83356 33236 83412 35756
rect 84476 35474 84532 35870
rect 84924 36484 84980 36494
rect 84924 35922 84980 36428
rect 84924 35870 84926 35922
rect 84978 35870 84980 35922
rect 84924 35812 84980 35870
rect 84924 35746 84980 35756
rect 86156 35812 86212 35822
rect 86156 35718 86212 35756
rect 86716 35810 86772 36540
rect 87052 36596 87108 36606
rect 87052 36502 87108 36540
rect 86716 35758 86718 35810
rect 86770 35758 86772 35810
rect 86716 35746 86772 35758
rect 87612 35810 87668 35822
rect 87612 35758 87614 35810
rect 87666 35758 87668 35810
rect 84476 35422 84478 35474
rect 84530 35422 84532 35474
rect 84476 35410 84532 35422
rect 85260 35474 85316 35486
rect 85260 35422 85262 35474
rect 85314 35422 85316 35474
rect 84252 34916 84308 34926
rect 84252 34822 84308 34860
rect 85260 34914 85316 35422
rect 85260 34862 85262 34914
rect 85314 34862 85316 34914
rect 85260 34850 85316 34862
rect 85596 35474 85652 35486
rect 85596 35422 85598 35474
rect 85650 35422 85652 35474
rect 85596 34916 85652 35422
rect 85596 34850 85652 34860
rect 85932 35474 85988 35486
rect 85932 35422 85934 35474
rect 85986 35422 85988 35474
rect 84476 34804 84532 34814
rect 84476 34710 84532 34748
rect 85148 34468 85204 34478
rect 83916 33908 83972 33918
rect 83916 33346 83972 33852
rect 83916 33294 83918 33346
rect 83970 33294 83972 33346
rect 83916 33282 83972 33294
rect 82908 33234 83412 33236
rect 82908 33182 82910 33234
rect 82962 33182 83412 33234
rect 82908 33180 83412 33182
rect 82908 32788 82964 33180
rect 83580 33124 83636 33134
rect 82908 32722 82964 32732
rect 83020 33122 83636 33124
rect 83020 33070 83582 33122
rect 83634 33070 83636 33122
rect 83020 33068 83636 33070
rect 83020 32674 83076 33068
rect 83580 33058 83636 33068
rect 84364 33122 84420 33134
rect 84364 33070 84366 33122
rect 84418 33070 84420 33122
rect 83020 32622 83022 32674
rect 83074 32622 83076 32674
rect 83020 32610 83076 32622
rect 83692 32788 83748 32798
rect 83132 30996 83188 31006
rect 83132 30902 83188 30940
rect 83692 29650 83748 32732
rect 84364 32788 84420 33070
rect 84364 32722 84420 32732
rect 85148 32450 85204 34412
rect 85932 34468 85988 35422
rect 86044 34804 86100 34814
rect 86044 34710 86100 34748
rect 85932 34402 85988 34412
rect 87500 34468 87556 34478
rect 86492 34244 86548 34254
rect 85820 34132 85876 34142
rect 85820 33346 85876 34076
rect 86492 33458 86548 34188
rect 86604 34132 86660 34142
rect 86604 34038 86660 34076
rect 86940 34132 86996 34142
rect 86492 33406 86494 33458
rect 86546 33406 86548 33458
rect 86492 33394 86548 33406
rect 86716 33684 86772 33694
rect 85820 33294 85822 33346
rect 85874 33294 85876 33346
rect 85820 33282 85876 33294
rect 85148 32398 85150 32450
rect 85202 32398 85204 32450
rect 85148 32386 85204 32398
rect 85596 33236 85652 33246
rect 85596 32786 85652 33180
rect 85596 32734 85598 32786
rect 85650 32734 85652 32786
rect 85596 32676 85652 32734
rect 86044 32788 86100 32798
rect 86044 32694 86100 32732
rect 86716 32786 86772 33628
rect 86716 32734 86718 32786
rect 86770 32734 86772 32786
rect 86716 32722 86772 32734
rect 84140 31666 84196 31678
rect 84140 31614 84142 31666
rect 84194 31614 84196 31666
rect 83804 31554 83860 31566
rect 83804 31502 83806 31554
rect 83858 31502 83860 31554
rect 83804 31108 83860 31502
rect 83916 31108 83972 31118
rect 83804 31106 83972 31108
rect 83804 31054 83918 31106
rect 83970 31054 83972 31106
rect 83804 31052 83972 31054
rect 83916 31042 83972 31052
rect 83692 29598 83694 29650
rect 83746 29598 83748 29650
rect 83692 29540 83748 29598
rect 84140 29652 84196 31614
rect 84588 30884 84644 30894
rect 84252 29652 84308 29662
rect 84140 29650 84308 29652
rect 84140 29598 84254 29650
rect 84306 29598 84308 29650
rect 84140 29596 84308 29598
rect 84252 29586 84308 29596
rect 83692 29474 83748 29484
rect 83244 29428 83300 29438
rect 83244 29334 83300 29372
rect 84588 29426 84644 30828
rect 85148 29540 85204 29550
rect 85148 29446 85204 29484
rect 84588 29374 84590 29426
rect 84642 29374 84644 29426
rect 84588 29362 84644 29374
rect 85372 29428 85428 29438
rect 85596 29428 85652 32620
rect 86940 31890 86996 34076
rect 87500 34020 87556 34412
rect 87612 34244 87668 35758
rect 87948 35812 88004 35822
rect 87612 34178 87668 34188
rect 87836 35698 87892 35710
rect 87836 35646 87838 35698
rect 87890 35646 87892 35698
rect 87612 34020 87668 34030
rect 87500 34018 87668 34020
rect 87500 33966 87614 34018
rect 87666 33966 87668 34018
rect 87500 33964 87668 33966
rect 87612 33954 87668 33964
rect 87276 33908 87332 33918
rect 87276 33814 87332 33852
rect 87836 33684 87892 35646
rect 87948 34242 88004 35756
rect 88060 34692 88116 47964
rect 88172 47684 88228 47694
rect 88172 47458 88228 47628
rect 88172 47406 88174 47458
rect 88226 47406 88228 47458
rect 88172 47394 88228 47406
rect 88396 46674 88452 48188
rect 88508 47236 88564 49868
rect 88620 48132 88676 48142
rect 88620 48038 88676 48076
rect 88508 47170 88564 47180
rect 88620 47346 88676 47358
rect 88620 47294 88622 47346
rect 88674 47294 88676 47346
rect 88396 46622 88398 46674
rect 88450 46622 88452 46674
rect 88396 46610 88452 46622
rect 88620 46004 88676 47294
rect 88620 45938 88676 45948
rect 88172 44994 88228 45006
rect 88172 44942 88174 44994
rect 88226 44942 88228 44994
rect 88172 41970 88228 44942
rect 88284 42532 88340 42542
rect 88284 42438 88340 42476
rect 88732 42530 88788 42542
rect 88732 42478 88734 42530
rect 88786 42478 88788 42530
rect 88732 42196 88788 42478
rect 88732 42130 88788 42140
rect 88172 41918 88174 41970
rect 88226 41918 88228 41970
rect 88172 40514 88228 41918
rect 88172 40462 88174 40514
rect 88226 40462 88228 40514
rect 88172 40292 88228 40462
rect 88172 40226 88228 40236
rect 88508 42084 88564 42094
rect 88508 39060 88564 42028
rect 88844 41300 88900 59724
rect 89404 59780 89460 59790
rect 89404 59686 89460 59724
rect 89628 59330 89684 59342
rect 89628 59278 89630 59330
rect 89682 59278 89684 59330
rect 89516 59218 89572 59230
rect 89516 59166 89518 59218
rect 89570 59166 89572 59218
rect 89292 58324 89348 58334
rect 89292 57538 89348 58268
rect 89292 57486 89294 57538
rect 89346 57486 89348 57538
rect 89292 57474 89348 57486
rect 89516 57204 89572 59166
rect 89516 57138 89572 57148
rect 89404 56866 89460 56878
rect 89404 56814 89406 56866
rect 89458 56814 89460 56866
rect 89068 55300 89124 55310
rect 89404 55300 89460 56814
rect 89628 56420 89684 59278
rect 89740 58996 89796 60508
rect 89852 59778 89908 59790
rect 89852 59726 89854 59778
rect 89906 59726 89908 59778
rect 89852 59444 89908 59726
rect 89852 59378 89908 59388
rect 89852 59220 89908 59230
rect 89852 59218 90132 59220
rect 89852 59166 89854 59218
rect 89906 59166 90132 59218
rect 89852 59164 90132 59166
rect 89852 59154 89908 59164
rect 89740 58940 90020 58996
rect 89628 56194 89684 56364
rect 89628 56142 89630 56194
rect 89682 56142 89684 56194
rect 89628 56130 89684 56142
rect 89740 56196 89796 56206
rect 89740 56194 89908 56196
rect 89740 56142 89742 56194
rect 89794 56142 89908 56194
rect 89740 56140 89908 56142
rect 89740 56130 89796 56140
rect 89740 55858 89796 55870
rect 89740 55806 89742 55858
rect 89794 55806 89796 55858
rect 89068 55298 89460 55300
rect 89068 55246 89070 55298
rect 89122 55246 89460 55298
rect 89068 55244 89460 55246
rect 89068 55234 89124 55244
rect 89292 54740 89348 54750
rect 89292 53058 89348 54684
rect 89404 53844 89460 55244
rect 89628 55748 89684 55758
rect 89516 54628 89572 54638
rect 89516 54534 89572 54572
rect 89628 54514 89684 55692
rect 89740 55410 89796 55806
rect 89740 55358 89742 55410
rect 89794 55358 89796 55410
rect 89740 55346 89796 55358
rect 89852 54740 89908 56140
rect 89852 54674 89908 54684
rect 89628 54462 89630 54514
rect 89682 54462 89684 54514
rect 89404 53778 89460 53788
rect 89516 54180 89572 54190
rect 89404 53172 89460 53182
rect 89516 53172 89572 54124
rect 89628 53844 89684 54462
rect 89964 54068 90020 58940
rect 90076 58548 90132 59164
rect 90076 58482 90132 58492
rect 90188 58996 90244 59006
rect 90076 56754 90132 56766
rect 90076 56702 90078 56754
rect 90130 56702 90132 56754
rect 90076 56308 90132 56702
rect 90076 56242 90132 56252
rect 90076 54514 90132 54526
rect 90076 54462 90078 54514
rect 90130 54462 90132 54514
rect 90076 54180 90132 54462
rect 90076 54114 90132 54124
rect 89964 54002 90020 54012
rect 89628 53788 90132 53844
rect 89964 53620 90020 53630
rect 89404 53170 89572 53172
rect 89404 53118 89406 53170
rect 89458 53118 89572 53170
rect 89404 53116 89572 53118
rect 89628 53618 90020 53620
rect 89628 53566 89966 53618
rect 90018 53566 90020 53618
rect 89628 53564 90020 53566
rect 89628 53170 89684 53564
rect 89964 53554 90020 53564
rect 89628 53118 89630 53170
rect 89682 53118 89684 53170
rect 89404 53106 89460 53116
rect 89628 53106 89684 53118
rect 89292 53006 89294 53058
rect 89346 53006 89348 53058
rect 89292 52994 89348 53006
rect 90076 52948 90132 53788
rect 90188 53060 90244 58940
rect 90300 56196 90356 56206
rect 90300 56102 90356 56140
rect 90412 55468 90468 63868
rect 90636 61010 90692 65548
rect 91196 64932 91252 67172
rect 91532 67170 91588 67790
rect 91756 67228 91812 72380
rect 91868 71652 91924 76412
rect 91980 75010 92036 75022
rect 91980 74958 91982 75010
rect 92034 74958 92036 75010
rect 91980 74340 92036 74958
rect 91980 74274 92036 74284
rect 92092 74788 92148 78932
rect 93212 78818 93268 78932
rect 93212 78766 93214 78818
rect 93266 78766 93268 78818
rect 93212 78754 93268 78766
rect 93548 78594 93604 78606
rect 93548 78542 93550 78594
rect 93602 78542 93604 78594
rect 93548 78146 93604 78542
rect 93548 78094 93550 78146
rect 93602 78094 93604 78146
rect 93548 78082 93604 78094
rect 93324 77250 93380 77262
rect 93324 77198 93326 77250
rect 93378 77198 93380 77250
rect 92540 77026 92596 77038
rect 92540 76974 92542 77026
rect 92594 76974 92596 77026
rect 92428 75794 92484 75806
rect 92428 75742 92430 75794
rect 92482 75742 92484 75794
rect 92316 75012 92372 75022
rect 92316 74918 92372 74956
rect 92092 74226 92148 74732
rect 92428 74676 92484 75742
rect 92428 74610 92484 74620
rect 92092 74174 92094 74226
rect 92146 74174 92148 74226
rect 92092 74162 92148 74174
rect 92540 74228 92596 76974
rect 93212 75794 93268 75806
rect 93212 75742 93214 75794
rect 93266 75742 93268 75794
rect 93212 75012 93268 75742
rect 93324 75124 93380 77198
rect 93548 77026 93604 77038
rect 93548 76974 93550 77026
rect 93602 76974 93604 77026
rect 93548 75796 93604 76974
rect 93548 75730 93604 75740
rect 93436 75124 93492 75134
rect 93324 75122 93492 75124
rect 93324 75070 93438 75122
rect 93490 75070 93492 75122
rect 93324 75068 93492 75070
rect 93436 75058 93492 75068
rect 93212 74946 93268 74956
rect 93772 74788 93828 78932
rect 94332 78932 94388 79326
rect 94332 78866 94388 78876
rect 94332 78034 94388 78046
rect 94332 77982 94334 78034
rect 94386 77982 94388 78034
rect 94332 77474 94388 77982
rect 94332 77422 94334 77474
rect 94386 77422 94388 77474
rect 94332 77410 94388 77422
rect 94444 78036 94500 80220
rect 94556 79714 94612 80668
rect 94556 79662 94558 79714
rect 94610 79662 94612 79714
rect 94556 79650 94612 79662
rect 94444 77364 94500 77980
rect 94668 77364 94724 77374
rect 94444 77362 94724 77364
rect 94444 77310 94670 77362
rect 94722 77310 94724 77362
rect 94444 77308 94724 77310
rect 94668 77298 94724 77308
rect 94444 77028 94500 77038
rect 93548 74676 93604 74686
rect 91868 71586 91924 71596
rect 91980 73442 92036 73454
rect 91980 73390 91982 73442
rect 92034 73390 92036 73442
rect 91980 71204 92036 73390
rect 91980 71138 92036 71148
rect 92316 73332 92372 73342
rect 92316 71202 92372 73276
rect 92540 72324 92596 74172
rect 93100 74340 93156 74350
rect 93100 74226 93156 74284
rect 93100 74174 93102 74226
rect 93154 74174 93156 74226
rect 93100 74162 93156 74174
rect 93548 74226 93604 74620
rect 93548 74174 93550 74226
rect 93602 74174 93604 74226
rect 93548 74162 93604 74174
rect 93772 74674 93828 74732
rect 93772 74622 93774 74674
rect 93826 74622 93828 74674
rect 93660 73444 93716 73454
rect 93660 73350 93716 73388
rect 92540 71876 92596 72268
rect 92316 71150 92318 71202
rect 92370 71150 92372 71202
rect 92316 71138 92372 71150
rect 92428 71874 92596 71876
rect 92428 71822 92542 71874
rect 92594 71822 92596 71874
rect 92428 71820 92596 71822
rect 91980 70980 92036 70990
rect 91980 70886 92036 70924
rect 92428 69410 92484 71820
rect 92540 71810 92596 71820
rect 92988 71204 93044 71214
rect 92988 70308 93044 71148
rect 93660 71092 93716 71102
rect 93660 70998 93716 71036
rect 93100 70980 93156 70990
rect 93100 70886 93156 70924
rect 93100 70308 93156 70318
rect 92988 70306 93156 70308
rect 92988 70254 93102 70306
rect 93154 70254 93156 70306
rect 92988 70252 93156 70254
rect 93100 70242 93156 70252
rect 92428 69358 92430 69410
rect 92482 69358 92484 69410
rect 92428 69346 92484 69358
rect 93436 69410 93492 69422
rect 93436 69358 93438 69410
rect 93490 69358 93492 69410
rect 93212 69300 93268 69310
rect 93212 69206 93268 69244
rect 93436 68964 93492 69358
rect 93436 68898 93492 68908
rect 91532 67118 91534 67170
rect 91586 67118 91588 67170
rect 91532 66276 91588 67118
rect 91532 66210 91588 66220
rect 91644 67172 91812 67228
rect 91868 68628 91924 68638
rect 91420 66164 91476 66202
rect 91420 66098 91476 66108
rect 91308 66052 91364 66062
rect 91308 65714 91364 65996
rect 91308 65662 91310 65714
rect 91362 65662 91364 65714
rect 91308 65650 91364 65662
rect 91196 64876 91364 64932
rect 90748 64820 90804 64830
rect 90748 64726 90804 64764
rect 91196 64482 91252 64494
rect 91196 64430 91198 64482
rect 91250 64430 91252 64482
rect 90748 63922 90804 63934
rect 90748 63870 90750 63922
rect 90802 63870 90804 63922
rect 90748 63700 90804 63870
rect 90748 62466 90804 63644
rect 90748 62414 90750 62466
rect 90802 62414 90804 62466
rect 90748 62402 90804 62414
rect 90860 63812 90916 63822
rect 90636 60958 90638 61010
rect 90690 60958 90692 61010
rect 90636 60946 90692 60958
rect 90636 58548 90692 58558
rect 90636 58454 90692 58492
rect 90524 56308 90580 56318
rect 90524 56214 90580 56252
rect 90636 56082 90692 56094
rect 90636 56030 90638 56082
rect 90690 56030 90692 56082
rect 90636 55748 90692 56030
rect 90636 55682 90692 55692
rect 90860 55468 90916 63756
rect 91196 63700 91252 64430
rect 91308 64148 91364 64876
rect 91308 63922 91364 64092
rect 91308 63870 91310 63922
rect 91362 63870 91364 63922
rect 91308 63858 91364 63870
rect 91196 63634 91252 63644
rect 91196 63140 91252 63150
rect 91196 63046 91252 63084
rect 91532 62354 91588 62366
rect 91532 62302 91534 62354
rect 91586 62302 91588 62354
rect 91532 62244 91588 62302
rect 91532 62178 91588 62188
rect 91644 61012 91700 67172
rect 91868 67060 91924 68572
rect 92092 68404 92148 68414
rect 92092 67954 92148 68348
rect 92092 67902 92094 67954
rect 92146 67902 92148 67954
rect 92092 67890 92148 67902
rect 93548 67956 93604 67966
rect 93548 67228 93604 67900
rect 91868 66386 91924 67004
rect 91868 66334 91870 66386
rect 91922 66334 91924 66386
rect 91868 65604 91924 66334
rect 93324 67172 93604 67228
rect 93212 66162 93268 66174
rect 93212 66110 93214 66162
rect 93266 66110 93268 66162
rect 91868 65538 91924 65548
rect 92540 66052 92596 66062
rect 93212 66052 93268 66110
rect 92540 66050 93268 66052
rect 92540 65998 92542 66050
rect 92594 65998 93268 66050
rect 92540 65996 93268 65998
rect 92316 63922 92372 63934
rect 92316 63870 92318 63922
rect 92370 63870 92372 63922
rect 92204 63252 92260 63262
rect 92204 63158 92260 63196
rect 91756 62916 91812 62926
rect 91756 62822 91812 62860
rect 92316 62916 92372 63870
rect 92540 63812 92596 65996
rect 92988 63924 93044 63934
rect 92988 63830 93044 63868
rect 92540 63746 92596 63756
rect 92316 62850 92372 62860
rect 93100 62468 93156 62478
rect 92316 62356 92372 62366
rect 92316 62262 92372 62300
rect 93100 62242 93156 62412
rect 93100 62190 93102 62242
rect 93154 62190 93156 62242
rect 92540 61460 92596 61470
rect 91644 60946 91700 60956
rect 91868 61236 91924 61246
rect 91756 59106 91812 59118
rect 91756 59054 91758 59106
rect 91810 59054 91812 59106
rect 91420 58436 91476 58446
rect 91420 58342 91476 58380
rect 91756 58436 91812 59054
rect 91756 58370 91812 58380
rect 91868 58212 91924 61180
rect 92428 60900 92484 60910
rect 92204 60564 92260 60574
rect 92204 60002 92260 60508
rect 92204 59950 92206 60002
rect 92258 59950 92260 60002
rect 92204 59938 92260 59950
rect 92316 59778 92372 59790
rect 92316 59726 92318 59778
rect 92370 59726 92372 59778
rect 91756 58156 91924 58212
rect 91980 58436 92036 58446
rect 91980 58210 92036 58380
rect 91980 58158 91982 58210
rect 92034 58158 92036 58210
rect 91420 57652 91476 57662
rect 91420 57558 91476 57596
rect 90412 55412 90692 55468
rect 90300 54628 90356 54638
rect 90300 54534 90356 54572
rect 90412 54516 90468 54526
rect 90188 52994 90244 53004
rect 90300 54068 90356 54078
rect 90076 52854 90132 52892
rect 90300 52724 90356 54012
rect 90412 53172 90468 54460
rect 90524 53172 90580 53182
rect 90412 53170 90580 53172
rect 90412 53118 90526 53170
rect 90578 53118 90580 53170
rect 90412 53116 90580 53118
rect 90524 53106 90580 53116
rect 90076 52668 90356 52724
rect 89180 52162 89236 52174
rect 89180 52110 89182 52162
rect 89234 52110 89236 52162
rect 89180 51156 89236 52110
rect 89852 52052 89908 52062
rect 90076 52052 90132 52668
rect 89852 52050 90132 52052
rect 89852 51998 89854 52050
rect 89906 51998 90132 52050
rect 89852 51996 90132 51998
rect 89852 51986 89908 51996
rect 89628 51940 89684 51950
rect 89628 51602 89684 51884
rect 89628 51550 89630 51602
rect 89682 51550 89684 51602
rect 89628 51538 89684 51550
rect 89964 51268 90020 51996
rect 89964 51174 90020 51212
rect 90188 51938 90244 51950
rect 90188 51886 90190 51938
rect 90242 51886 90244 51938
rect 90188 51828 90244 51886
rect 89516 51156 89572 51166
rect 89180 51154 89572 51156
rect 89180 51102 89518 51154
rect 89570 51102 89572 51154
rect 89180 51100 89572 51102
rect 88956 50482 89012 50494
rect 88956 50430 88958 50482
rect 89010 50430 89012 50482
rect 88956 49812 89012 50430
rect 88956 49746 89012 49756
rect 89068 50484 89124 50494
rect 89068 49140 89124 50428
rect 89068 49074 89124 49084
rect 89068 46004 89124 46014
rect 89068 45910 89124 45948
rect 88396 39058 88564 39060
rect 88396 39006 88510 39058
rect 88562 39006 88564 39058
rect 88396 39004 88564 39006
rect 88172 36596 88228 36606
rect 88172 35026 88228 36540
rect 88172 34974 88174 35026
rect 88226 34974 88228 35026
rect 88172 34962 88228 34974
rect 88060 34626 88116 34636
rect 87948 34190 87950 34242
rect 88002 34190 88004 34242
rect 87948 34178 88004 34190
rect 88172 34242 88228 34254
rect 88172 34190 88174 34242
rect 88226 34190 88228 34242
rect 87836 33618 87892 33628
rect 88172 32788 88228 34190
rect 88396 34132 88452 39004
rect 88508 38994 88564 39004
rect 88732 41244 88900 41300
rect 88508 37828 88564 37838
rect 88508 37734 88564 37772
rect 88732 36596 88788 41244
rect 88844 41074 88900 41086
rect 88844 41022 88846 41074
rect 88898 41022 88900 41074
rect 88844 40628 88900 41022
rect 88844 40562 88900 40572
rect 89180 38276 89236 51100
rect 89516 51090 89572 51100
rect 90188 51044 90244 51772
rect 90412 51266 90468 51278
rect 90412 51214 90414 51266
rect 90466 51214 90468 51266
rect 90412 51154 90468 51214
rect 90412 51102 90414 51154
rect 90466 51102 90468 51154
rect 90412 51090 90468 51102
rect 89964 50988 90244 51044
rect 89292 50484 89348 50494
rect 89292 50390 89348 50428
rect 89964 50482 90020 50988
rect 89964 50430 89966 50482
rect 90018 50430 90020 50482
rect 89964 50418 90020 50430
rect 90076 50708 90132 50718
rect 90076 50482 90132 50652
rect 90076 50430 90078 50482
rect 90130 50430 90132 50482
rect 89740 50372 89796 50382
rect 89404 50370 89796 50372
rect 89404 50318 89742 50370
rect 89794 50318 89796 50370
rect 89404 50316 89796 50318
rect 89404 50034 89460 50316
rect 89740 50306 89796 50316
rect 90076 50372 90132 50430
rect 90076 50306 90132 50316
rect 90188 50484 90244 50494
rect 89404 49982 89406 50034
rect 89458 49982 89460 50034
rect 89404 49970 89460 49982
rect 90188 50034 90244 50428
rect 90188 49982 90190 50034
rect 90242 49982 90244 50034
rect 90188 49970 90244 49982
rect 90300 49924 90356 49934
rect 90300 49830 90356 49868
rect 89292 49812 89348 49822
rect 89292 48804 89348 49756
rect 89628 49812 89684 49822
rect 89628 49810 90132 49812
rect 89628 49758 89630 49810
rect 89682 49758 90132 49810
rect 89628 49756 90132 49758
rect 89628 49746 89684 49756
rect 89292 48738 89348 48748
rect 90076 48354 90132 49756
rect 90076 48302 90078 48354
rect 90130 48302 90132 48354
rect 90076 48290 90132 48302
rect 90188 49586 90244 49598
rect 90188 49534 90190 49586
rect 90242 49534 90244 49586
rect 89292 48242 89348 48254
rect 89292 48190 89294 48242
rect 89346 48190 89348 48242
rect 89292 47458 89348 48190
rect 89964 47572 90020 47582
rect 90188 47572 90244 49534
rect 89964 47570 90244 47572
rect 89964 47518 89966 47570
rect 90018 47518 90244 47570
rect 89964 47516 90244 47518
rect 89964 47506 90020 47516
rect 89292 47406 89294 47458
rect 89346 47406 89348 47458
rect 89292 46676 89348 47406
rect 89740 47236 89796 47246
rect 89628 46676 89684 46686
rect 89292 46674 89684 46676
rect 89292 46622 89630 46674
rect 89682 46622 89684 46674
rect 89292 46620 89684 46622
rect 89628 45668 89684 46620
rect 89740 45892 89796 47180
rect 89740 45760 89796 45836
rect 89852 47124 89908 47134
rect 89852 45778 89908 47068
rect 90412 46564 90468 46574
rect 90076 46562 90468 46564
rect 90076 46510 90414 46562
rect 90466 46510 90468 46562
rect 90076 46508 90468 46510
rect 90076 45890 90132 46508
rect 90412 46498 90468 46508
rect 90636 46340 90692 55412
rect 90748 55412 90916 55468
rect 90748 54068 90804 55412
rect 90860 54740 90916 54750
rect 90860 54646 90916 54684
rect 91084 54628 91140 54638
rect 91084 54534 91140 54572
rect 91196 54516 91252 54526
rect 91252 54460 91364 54516
rect 91196 54384 91252 54460
rect 90748 54012 90916 54068
rect 90748 53844 90804 53854
rect 90748 53730 90804 53788
rect 90748 53678 90750 53730
rect 90802 53678 90804 53730
rect 90748 53666 90804 53678
rect 90860 53732 90916 54012
rect 90860 52834 90916 53676
rect 91196 53844 91252 53854
rect 91308 53844 91364 54460
rect 91644 54402 91700 54414
rect 91644 54350 91646 54402
rect 91698 54350 91700 54402
rect 91644 54292 91700 54350
rect 91644 54226 91700 54236
rect 91644 53844 91700 53854
rect 91308 53842 91700 53844
rect 91308 53790 91646 53842
rect 91698 53790 91700 53842
rect 91308 53788 91700 53790
rect 91196 53730 91252 53788
rect 91644 53778 91700 53788
rect 91196 53678 91198 53730
rect 91250 53678 91252 53730
rect 91196 53666 91252 53678
rect 90860 52782 90862 52834
rect 90914 52782 90916 52834
rect 90860 52164 90916 52782
rect 91196 52164 91252 52174
rect 90860 52162 91364 52164
rect 90860 52110 91198 52162
rect 91250 52110 91364 52162
rect 90860 52108 91364 52110
rect 91196 52098 91252 52108
rect 91084 50596 91140 50606
rect 91084 50502 91140 50540
rect 90748 50370 90804 50382
rect 90748 50318 90750 50370
rect 90802 50318 90804 50370
rect 90748 49924 90804 50318
rect 90748 49858 90804 49868
rect 90972 50370 91028 50382
rect 90972 50318 90974 50370
rect 91026 50318 91028 50370
rect 90972 47572 91028 50318
rect 91196 50372 91252 50382
rect 91196 50036 91252 50316
rect 91308 50260 91364 52108
rect 91756 52052 91812 58156
rect 91980 57652 92036 58158
rect 92316 57764 92372 59726
rect 92428 58436 92484 60844
rect 92540 60002 92596 61404
rect 92540 59950 92542 60002
rect 92594 59950 92596 60002
rect 92540 59938 92596 59950
rect 93100 58436 93156 62190
rect 93212 62244 93268 62254
rect 93212 61684 93268 62188
rect 93212 61590 93268 61628
rect 93324 61236 93380 67172
rect 93772 66948 93828 74622
rect 93996 75010 94052 75022
rect 93996 74958 93998 75010
rect 94050 74958 94052 75010
rect 93996 74004 94052 74958
rect 94332 75012 94388 75022
rect 94332 74918 94388 74956
rect 93996 73890 94052 73948
rect 93996 73838 93998 73890
rect 94050 73838 94052 73890
rect 93996 73444 94052 73838
rect 93996 73378 94052 73388
rect 94220 73218 94276 73230
rect 94220 73166 94222 73218
rect 94274 73166 94276 73218
rect 94220 73106 94276 73166
rect 94220 73054 94222 73106
rect 94274 73054 94276 73106
rect 94220 73042 94276 73054
rect 94108 72324 94164 72334
rect 93996 71092 94052 71102
rect 94108 71092 94164 72268
rect 93884 71090 94164 71092
rect 93884 71038 93998 71090
rect 94050 71038 94164 71090
rect 93884 71036 94164 71038
rect 93884 70196 93940 71036
rect 93996 71026 94052 71036
rect 93884 70194 94164 70196
rect 93884 70142 93886 70194
rect 93938 70142 94164 70194
rect 93884 70140 94164 70142
rect 93884 70130 93940 70140
rect 94108 69522 94164 70140
rect 94108 69470 94110 69522
rect 94162 69470 94164 69522
rect 94108 69458 94164 69470
rect 93996 67060 94052 67070
rect 93996 66966 94052 67004
rect 93548 66892 93772 66948
rect 93548 66162 93604 66892
rect 93772 66882 93828 66892
rect 94108 66836 94164 66846
rect 94108 66388 94164 66780
rect 94108 66294 94164 66332
rect 93548 66110 93550 66162
rect 93602 66110 93604 66162
rect 93548 66098 93604 66110
rect 94332 65492 94388 65502
rect 94332 65398 94388 65436
rect 93772 65378 93828 65390
rect 93772 65326 93774 65378
rect 93826 65326 93828 65378
rect 93772 65044 93828 65326
rect 93772 64978 93828 64988
rect 94220 65044 94276 65054
rect 94220 64818 94276 64988
rect 94220 64766 94222 64818
rect 94274 64766 94276 64818
rect 94220 64754 94276 64766
rect 93660 64484 93716 64494
rect 93660 64390 93716 64428
rect 94444 64484 94500 76972
rect 94780 77028 94836 81004
rect 94892 80388 94948 82574
rect 95116 82180 95172 86492
rect 95564 86482 95620 86492
rect 95900 86436 95956 86446
rect 95900 86434 96068 86436
rect 95900 86382 95902 86434
rect 95954 86382 96068 86434
rect 95900 86380 96068 86382
rect 95900 86370 95956 86380
rect 95900 85988 95956 85998
rect 95676 85986 95956 85988
rect 95676 85934 95902 85986
rect 95954 85934 95956 85986
rect 95676 85932 95956 85934
rect 95564 85876 95620 85886
rect 95228 85874 95620 85876
rect 95228 85822 95566 85874
rect 95618 85822 95620 85874
rect 95228 85820 95620 85822
rect 95228 84530 95284 85820
rect 95564 85810 95620 85820
rect 95676 85202 95732 85932
rect 95900 85922 95956 85932
rect 95676 85150 95678 85202
rect 95730 85150 95732 85202
rect 95676 85138 95732 85150
rect 96012 84980 96068 86380
rect 96636 85484 96900 85494
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96636 85418 96900 85428
rect 95676 84924 96068 84980
rect 95228 84478 95230 84530
rect 95282 84478 95284 84530
rect 95228 84466 95284 84478
rect 95564 84532 95620 84542
rect 95564 84306 95620 84476
rect 95564 84254 95566 84306
rect 95618 84254 95620 84306
rect 95564 84242 95620 84254
rect 95676 83634 95732 84924
rect 95676 83582 95678 83634
rect 95730 83582 95732 83634
rect 95676 83570 95732 83582
rect 95788 84418 95844 84430
rect 95788 84366 95790 84418
rect 95842 84366 95844 84418
rect 95788 83636 95844 84366
rect 95228 82180 95284 82190
rect 95116 82178 95284 82180
rect 95116 82126 95230 82178
rect 95282 82126 95284 82178
rect 95116 82124 95284 82126
rect 95228 82114 95284 82124
rect 95788 82180 95844 83580
rect 96348 84420 96404 84430
rect 95564 81954 95620 81966
rect 95564 81902 95566 81954
rect 95618 81902 95620 81954
rect 95564 81844 95620 81902
rect 95340 81788 95620 81844
rect 94892 80294 94948 80332
rect 95228 80946 95284 80958
rect 95228 80894 95230 80946
rect 95282 80894 95284 80946
rect 94892 79716 94948 79726
rect 94892 79622 94948 79660
rect 95228 79716 95284 80894
rect 95340 80500 95396 81788
rect 95788 81282 95844 82124
rect 96236 83524 96292 83534
rect 96236 81954 96292 83468
rect 96236 81902 96238 81954
rect 96290 81902 96292 81954
rect 96236 81620 96292 81902
rect 96348 81842 96404 84364
rect 96636 83916 96900 83926
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96636 83850 96900 83860
rect 96636 82348 96900 82358
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96636 82282 96900 82292
rect 97356 82068 97412 82078
rect 97356 81974 97412 82012
rect 96348 81790 96350 81842
rect 96402 81790 96404 81842
rect 96348 81778 96404 81790
rect 96908 81730 96964 81742
rect 96908 81678 96910 81730
rect 96962 81678 96964 81730
rect 96908 81620 96964 81678
rect 96236 81564 96964 81620
rect 95788 81230 95790 81282
rect 95842 81230 95844 81282
rect 95564 81060 95620 81070
rect 95340 79940 95396 80444
rect 95340 79874 95396 79884
rect 95452 80612 95508 80622
rect 95228 79650 95284 79660
rect 94780 76962 94836 76972
rect 94892 78818 94948 78830
rect 94892 78766 94894 78818
rect 94946 78766 94948 78818
rect 94892 77474 94948 78766
rect 95452 78146 95508 80556
rect 95564 78596 95620 81004
rect 95676 80274 95732 80286
rect 95676 80222 95678 80274
rect 95730 80222 95732 80274
rect 95676 79828 95732 80222
rect 95788 80276 95844 81230
rect 96124 81282 96180 81294
rect 96124 81230 96126 81282
rect 96178 81230 96180 81282
rect 96124 80612 96180 81230
rect 97244 81060 97300 81070
rect 97244 80966 97300 81004
rect 96636 80780 96900 80790
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96636 80714 96900 80724
rect 96124 80546 96180 80556
rect 95788 80210 95844 80220
rect 95676 79762 95732 79772
rect 97244 79828 97300 79838
rect 97244 79734 97300 79772
rect 95788 79714 95844 79726
rect 95788 79662 95790 79714
rect 95842 79662 95844 79714
rect 95788 78988 95844 79662
rect 96124 79716 96180 79726
rect 96124 79622 96180 79660
rect 95676 78932 95844 78988
rect 96348 79604 96404 79614
rect 95676 78930 95732 78932
rect 95676 78878 95678 78930
rect 95730 78878 95732 78930
rect 95676 78866 95732 78878
rect 95564 78530 95620 78540
rect 96348 78258 96404 79548
rect 96636 79212 96900 79222
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96636 79146 96900 79156
rect 96348 78206 96350 78258
rect 96402 78206 96404 78258
rect 96348 78194 96404 78206
rect 95452 78094 95454 78146
rect 95506 78094 95508 78146
rect 95452 78082 95508 78094
rect 95228 78036 95284 78046
rect 95228 77942 95284 77980
rect 94892 77422 94894 77474
rect 94946 77422 94948 77474
rect 94892 76354 94948 77422
rect 96012 77810 96068 77822
rect 96012 77758 96014 77810
rect 96066 77758 96068 77810
rect 95004 77028 95060 77038
rect 95004 76934 95060 76972
rect 96012 77028 96068 77758
rect 96636 77644 96900 77654
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96636 77578 96900 77588
rect 96012 76962 96068 76972
rect 97132 77028 97188 77038
rect 94892 76302 94894 76354
rect 94946 76302 94948 76354
rect 94892 75684 94948 76302
rect 97132 76354 97188 76972
rect 97132 76302 97134 76354
rect 97186 76302 97188 76354
rect 96636 76076 96900 76086
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96636 76010 96900 76020
rect 97132 75906 97188 76302
rect 97132 75854 97134 75906
rect 97186 75854 97188 75906
rect 97132 75842 97188 75854
rect 95340 75796 95396 75806
rect 95340 75702 95396 75740
rect 94556 75012 94612 75022
rect 94556 72436 94612 74956
rect 94892 74114 94948 75628
rect 96012 75684 96068 75694
rect 96012 75590 96068 75628
rect 97356 75570 97412 75582
rect 97356 75518 97358 75570
rect 97410 75518 97412 75570
rect 96796 75460 96852 75470
rect 95900 75458 96852 75460
rect 95900 75406 96798 75458
rect 96850 75406 96852 75458
rect 95900 75404 96852 75406
rect 95564 75010 95620 75022
rect 95564 74958 95566 75010
rect 95618 74958 95620 75010
rect 95564 74228 95620 74958
rect 95900 75010 95956 75404
rect 96796 75394 96852 75404
rect 95900 74958 95902 75010
rect 95954 74958 95956 75010
rect 95900 74946 95956 74958
rect 96348 74788 96404 74798
rect 96348 74694 96404 74732
rect 97132 74788 97188 74798
rect 97356 74788 97412 75518
rect 97132 74786 97412 74788
rect 97132 74734 97134 74786
rect 97186 74734 97412 74786
rect 97132 74732 97412 74734
rect 96636 74508 96900 74518
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96636 74442 96900 74452
rect 95676 74228 95732 74238
rect 95564 74226 95732 74228
rect 95564 74174 95678 74226
rect 95730 74174 95732 74226
rect 95564 74172 95732 74174
rect 95676 74162 95732 74172
rect 96348 74228 96404 74238
rect 94892 74062 94894 74114
rect 94946 74062 94948 74114
rect 94892 74050 94948 74062
rect 95788 74004 95844 74014
rect 95788 73442 95844 73948
rect 95788 73390 95790 73442
rect 95842 73390 95844 73442
rect 95788 73378 95844 73390
rect 96348 73442 96404 74172
rect 97132 74004 97188 74732
rect 97132 73938 97188 73948
rect 97244 73444 97300 73454
rect 96348 73390 96350 73442
rect 96402 73390 96404 73442
rect 96348 73378 96404 73390
rect 97020 73442 97300 73444
rect 97020 73390 97246 73442
rect 97298 73390 97300 73442
rect 97020 73388 97300 73390
rect 95228 73332 95284 73342
rect 95228 73238 95284 73276
rect 94668 73218 94724 73230
rect 94668 73166 94670 73218
rect 94722 73166 94724 73218
rect 94668 72548 94724 73166
rect 94668 72482 94724 72492
rect 94892 73106 94948 73118
rect 94892 73054 94894 73106
rect 94946 73054 94948 73106
rect 94892 72660 94948 73054
rect 95564 73106 95620 73118
rect 95564 73054 95566 73106
rect 95618 73054 95620 73106
rect 95564 72660 95620 73054
rect 96636 72940 96900 72950
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96636 72874 96900 72884
rect 94892 72658 95620 72660
rect 94892 72606 94894 72658
rect 94946 72606 95620 72658
rect 94892 72604 95620 72606
rect 97020 72658 97076 73388
rect 97244 73378 97300 73388
rect 97020 72606 97022 72658
rect 97074 72606 97076 72658
rect 94556 72370 94612 72380
rect 94780 70866 94836 70878
rect 94780 70814 94782 70866
rect 94834 70814 94836 70866
rect 94780 70418 94836 70814
rect 94780 70366 94782 70418
rect 94834 70366 94836 70418
rect 94780 70354 94836 70366
rect 94892 70196 94948 72604
rect 97020 72594 97076 72606
rect 95564 71652 95620 71662
rect 95564 71558 95620 71596
rect 96636 71372 96900 71382
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96636 71306 96900 71316
rect 95004 71092 95060 71102
rect 95004 70308 95060 71036
rect 96460 71092 96516 71102
rect 96460 70998 96516 71036
rect 95116 70868 95172 70878
rect 95116 70866 95620 70868
rect 95116 70814 95118 70866
rect 95170 70814 95620 70866
rect 95116 70812 95620 70814
rect 95116 70802 95172 70812
rect 95340 70308 95396 70318
rect 95004 70306 95396 70308
rect 95004 70254 95342 70306
rect 95394 70254 95396 70306
rect 95004 70252 95396 70254
rect 95340 70242 95396 70252
rect 95452 70308 95508 70318
rect 94892 70140 95060 70196
rect 94892 69524 94948 69534
rect 94892 69430 94948 69468
rect 94668 67844 94724 67854
rect 94668 66274 94724 67788
rect 95004 67228 95060 70140
rect 95116 70084 95172 70094
rect 95116 67956 95172 70028
rect 95116 67890 95172 67900
rect 95340 69524 95396 69534
rect 95004 67172 95172 67228
rect 95116 66388 95172 67172
rect 95340 67170 95396 69468
rect 95340 67118 95342 67170
rect 95394 67118 95396 67170
rect 95340 67106 95396 67118
rect 95452 67172 95508 70252
rect 95564 67956 95620 70812
rect 95676 70866 95732 70878
rect 95676 70814 95678 70866
rect 95730 70814 95732 70866
rect 95676 70532 95732 70814
rect 95676 70466 95732 70476
rect 96012 70754 96068 70766
rect 96012 70702 96014 70754
rect 96066 70702 96068 70754
rect 95676 70306 95732 70318
rect 95676 70254 95678 70306
rect 95730 70254 95732 70306
rect 95676 69524 95732 70254
rect 95676 69458 95732 69468
rect 96012 69524 96068 70702
rect 96460 70196 96516 70206
rect 96012 69458 96068 69468
rect 96236 70140 96460 70196
rect 96236 68738 96292 70140
rect 96460 70102 96516 70140
rect 97132 70084 97188 70094
rect 97132 69990 97188 70028
rect 96636 69804 96900 69814
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96636 69738 96900 69748
rect 97020 69524 97076 69534
rect 97020 69430 97076 69468
rect 96236 68686 96238 68738
rect 96290 68686 96292 68738
rect 95676 67956 95732 67966
rect 95564 67954 95732 67956
rect 95564 67902 95678 67954
rect 95730 67902 95732 67954
rect 95564 67900 95732 67902
rect 95676 67890 95732 67900
rect 96236 67844 96292 68686
rect 96636 68236 96900 68246
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96636 68170 96900 68180
rect 96348 67844 96404 67854
rect 96236 67788 96348 67844
rect 96348 67712 96404 67788
rect 97356 67844 97412 67854
rect 97356 67750 97412 67788
rect 96908 67618 96964 67630
rect 96908 67566 96910 67618
rect 96962 67566 96964 67618
rect 95452 67106 95508 67116
rect 96348 67172 96404 67182
rect 96348 67078 96404 67116
rect 95228 67058 95284 67070
rect 95228 67006 95230 67058
rect 95282 67006 95284 67058
rect 95228 66836 95284 67006
rect 95228 66770 95284 66780
rect 95788 67060 95844 67070
rect 95116 66332 95620 66388
rect 94668 66222 94670 66274
rect 94722 66222 94724 66274
rect 94668 66210 94724 66222
rect 95452 66164 95508 66174
rect 94780 66162 95508 66164
rect 94780 66110 95454 66162
rect 95506 66110 95508 66162
rect 94780 66108 95508 66110
rect 94780 65828 94836 66108
rect 95452 66098 95508 66108
rect 94556 65772 94836 65828
rect 94556 65714 94612 65772
rect 94556 65662 94558 65714
rect 94610 65662 94612 65714
rect 94556 65650 94612 65662
rect 95340 65492 95396 65502
rect 95564 65492 95620 66332
rect 94444 64418 94500 64428
rect 95228 65266 95284 65278
rect 95228 65214 95230 65266
rect 95282 65214 95284 65266
rect 93436 64148 93492 64158
rect 93436 64054 93492 64092
rect 94556 64148 94612 64158
rect 94556 64054 94612 64092
rect 94332 63924 94388 63934
rect 95228 63924 95284 65214
rect 94332 63922 95284 63924
rect 94332 63870 94334 63922
rect 94386 63870 95284 63922
rect 94332 63868 95284 63870
rect 94332 63858 94388 63868
rect 95228 63700 95284 63710
rect 95340 63700 95396 65436
rect 95228 63698 95396 63700
rect 95228 63646 95230 63698
rect 95282 63646 95396 63698
rect 95228 63644 95396 63646
rect 95452 65436 95620 65492
rect 95228 63634 95284 63644
rect 95004 63140 95060 63150
rect 94332 63026 94388 63038
rect 94332 62974 94334 63026
rect 94386 62974 94388 63026
rect 93660 62914 93716 62926
rect 93660 62862 93662 62914
rect 93714 62862 93716 62914
rect 93660 62692 93716 62862
rect 93996 62916 94052 62926
rect 94220 62916 94276 62926
rect 93996 62914 94164 62916
rect 93996 62862 93998 62914
rect 94050 62862 94164 62914
rect 93996 62860 94164 62862
rect 93996 62850 94052 62860
rect 93660 62626 93716 62636
rect 93660 62354 93716 62366
rect 93660 62302 93662 62354
rect 93714 62302 93716 62354
rect 93660 61572 93716 62302
rect 93884 61572 93940 61582
rect 93660 61570 93940 61572
rect 93660 61518 93886 61570
rect 93938 61518 93940 61570
rect 93660 61516 93940 61518
rect 93324 61170 93380 61180
rect 93548 60676 93604 60686
rect 93884 60676 93940 61516
rect 93548 60674 93940 60676
rect 93548 60622 93550 60674
rect 93602 60622 93940 60674
rect 93548 60620 93940 60622
rect 93548 60002 93604 60620
rect 94108 60564 94164 62860
rect 94220 62822 94276 62860
rect 94332 62692 94388 62974
rect 95004 63026 95060 63084
rect 95004 62974 95006 63026
rect 95058 62974 95060 63026
rect 95004 62962 95060 62974
rect 95116 63026 95172 63038
rect 95116 62974 95118 63026
rect 95170 62974 95172 63026
rect 94780 62916 94836 62926
rect 94332 62626 94388 62636
rect 94556 62914 94836 62916
rect 94556 62862 94782 62914
rect 94834 62862 94836 62914
rect 94556 62860 94836 62862
rect 94332 62244 94388 62254
rect 94108 60498 94164 60508
rect 94220 62242 94388 62244
rect 94220 62190 94334 62242
rect 94386 62190 94388 62242
rect 94220 62188 94388 62190
rect 93548 59950 93550 60002
rect 93602 59950 93604 60002
rect 93548 59938 93604 59950
rect 94220 59442 94276 62188
rect 94332 62178 94388 62188
rect 94332 60004 94388 60014
rect 94332 59910 94388 59948
rect 94220 59390 94222 59442
rect 94274 59390 94276 59442
rect 94220 59378 94276 59390
rect 94444 59332 94500 59342
rect 94444 59238 94500 59276
rect 94556 59330 94612 62860
rect 94780 62850 94836 62860
rect 95116 62692 95172 62974
rect 95116 62626 95172 62636
rect 95452 61684 95508 65436
rect 95564 65266 95620 65278
rect 95564 65214 95566 65266
rect 95618 65214 95620 65266
rect 95564 65044 95620 65214
rect 95564 64978 95620 64988
rect 95452 61618 95508 61628
rect 95564 64484 95620 64494
rect 95564 63698 95620 64428
rect 95564 63646 95566 63698
rect 95618 63646 95620 63698
rect 94668 61460 94724 61470
rect 95564 61460 95620 63646
rect 95676 62914 95732 62926
rect 95676 62862 95678 62914
rect 95730 62862 95732 62914
rect 95676 62692 95732 62862
rect 95676 62626 95732 62636
rect 94668 61366 94724 61404
rect 95452 61404 95620 61460
rect 94556 59278 94558 59330
rect 94610 59278 94612 59330
rect 94556 59266 94612 59278
rect 92428 58380 92596 58436
rect 92316 57698 92372 57708
rect 92428 58210 92484 58222
rect 92428 58158 92430 58210
rect 92482 58158 92484 58210
rect 92204 57652 92260 57662
rect 91980 57596 92204 57652
rect 92204 57558 92260 57596
rect 92428 57652 92484 58158
rect 92428 57586 92484 57596
rect 92204 56978 92260 56990
rect 92204 56926 92206 56978
rect 92258 56926 92260 56978
rect 91868 56644 91924 56654
rect 91868 55410 91924 56588
rect 92204 56308 92260 56926
rect 92204 56242 92260 56252
rect 92316 56082 92372 56094
rect 92316 56030 92318 56082
rect 92370 56030 92372 56082
rect 91868 55358 91870 55410
rect 91922 55358 91924 55410
rect 91868 55346 91924 55358
rect 91980 55972 92036 55982
rect 91756 51986 91812 51996
rect 91868 53956 91924 53966
rect 91420 51938 91476 51950
rect 91420 51886 91422 51938
rect 91474 51886 91476 51938
rect 91420 51828 91476 51886
rect 91868 51938 91924 53900
rect 91868 51886 91870 51938
rect 91922 51886 91924 51938
rect 91868 51828 91924 51886
rect 91420 51772 91924 51828
rect 91532 50484 91588 50494
rect 91532 50390 91588 50428
rect 91756 50370 91812 51772
rect 91980 51378 92036 55916
rect 92316 55972 92372 56030
rect 92316 55906 92372 55916
rect 92316 55748 92372 55758
rect 92316 55410 92372 55692
rect 92316 55358 92318 55410
rect 92370 55358 92372 55410
rect 92316 55346 92372 55358
rect 92204 55300 92260 55310
rect 92092 54404 92148 54414
rect 92092 53956 92148 54348
rect 92092 53890 92148 53900
rect 92204 53844 92260 55244
rect 92204 53170 92260 53788
rect 92316 54852 92372 54862
rect 92316 53730 92372 54796
rect 92316 53678 92318 53730
rect 92370 53678 92372 53730
rect 92316 53666 92372 53678
rect 92540 53732 92596 58380
rect 92204 53118 92206 53170
rect 92258 53118 92260 53170
rect 92204 53106 92260 53118
rect 92540 52836 92596 53676
rect 92652 58380 93156 58436
rect 92652 53060 92708 58380
rect 94892 58324 94948 58334
rect 94892 58230 94948 58268
rect 93212 58212 93268 58222
rect 93212 58210 93492 58212
rect 93212 58158 93214 58210
rect 93266 58158 93492 58210
rect 93212 58156 93492 58158
rect 93212 58146 93268 58156
rect 92764 57764 92820 57774
rect 92764 57670 92820 57708
rect 92876 57764 92932 57774
rect 92876 57762 93044 57764
rect 92876 57710 92878 57762
rect 92930 57710 93044 57762
rect 92876 57708 93044 57710
rect 92876 57698 92932 57708
rect 92764 54852 92820 54862
rect 92764 54626 92820 54796
rect 92988 54740 93044 57708
rect 93100 57650 93156 57662
rect 93100 57598 93102 57650
rect 93154 57598 93156 57650
rect 93100 56980 93156 57598
rect 93100 56914 93156 56924
rect 93436 56866 93492 58156
rect 94556 58210 94612 58222
rect 94556 58158 94558 58210
rect 94610 58158 94612 58210
rect 94332 57764 94388 57774
rect 94332 57670 94388 57708
rect 93436 56814 93438 56866
rect 93490 56814 93492 56866
rect 93100 56642 93156 56654
rect 93100 56590 93102 56642
rect 93154 56590 93156 56642
rect 93100 56420 93156 56590
rect 93324 56644 93380 56654
rect 93324 56550 93380 56588
rect 93100 56354 93156 56364
rect 93436 55748 93492 56814
rect 93660 57652 93716 57662
rect 93660 56868 93716 57596
rect 93660 56802 93716 56812
rect 94332 56868 94388 56878
rect 93884 56644 93940 56654
rect 93436 55682 93492 55692
rect 93548 55860 93604 55870
rect 93548 55300 93604 55804
rect 93548 55168 93604 55244
rect 93548 54852 93604 54862
rect 93100 54740 93156 54750
rect 92988 54738 93156 54740
rect 92988 54686 93102 54738
rect 93154 54686 93156 54738
rect 92988 54684 93156 54686
rect 93100 54674 93156 54684
rect 92764 54574 92766 54626
rect 92818 54574 92820 54626
rect 92764 54562 92820 54574
rect 92876 54626 92932 54638
rect 92876 54574 92878 54626
rect 92930 54574 92932 54626
rect 92876 53956 92932 54574
rect 93548 54626 93604 54796
rect 93884 54738 93940 56588
rect 94332 55860 94388 56812
rect 94332 55794 94388 55804
rect 94556 55468 94612 58158
rect 94332 55412 94388 55422
rect 94444 55412 94612 55468
rect 94780 58210 94836 58222
rect 94780 58158 94782 58210
rect 94834 58158 94836 58210
rect 94332 55410 94500 55412
rect 94332 55358 94334 55410
rect 94386 55358 94500 55410
rect 94332 55356 94500 55358
rect 94332 55346 94388 55356
rect 93884 54686 93886 54738
rect 93938 54686 93940 54738
rect 93884 54674 93940 54686
rect 94668 54740 94724 54750
rect 94780 54740 94836 58158
rect 95340 58210 95396 58222
rect 95340 58158 95342 58210
rect 95394 58158 95396 58210
rect 95340 57764 95396 58158
rect 95340 57698 95396 57708
rect 95004 56980 95060 56990
rect 95004 56886 95060 56924
rect 95452 55468 95508 61404
rect 95788 60786 95844 67004
rect 96908 67060 96964 67566
rect 96908 66994 96964 67004
rect 96012 66948 96068 66958
rect 96012 66854 96068 66892
rect 97132 66948 97188 66958
rect 97132 66854 97188 66892
rect 96124 66836 96180 66846
rect 96124 65492 96180 66780
rect 96636 66668 96900 66678
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96636 66602 96900 66612
rect 97468 66500 97524 96012
rect 97804 85202 97860 85214
rect 97804 85150 97806 85202
rect 97858 85150 97860 85202
rect 97804 84420 97860 85150
rect 97804 84354 97860 84364
rect 97804 83634 97860 83646
rect 97804 83582 97806 83634
rect 97858 83582 97860 83634
rect 97804 81732 97860 83582
rect 97692 81730 97860 81732
rect 97692 81678 97806 81730
rect 97858 81678 97860 81730
rect 97692 81676 97860 81678
rect 97692 80500 97748 81676
rect 97804 81666 97860 81676
rect 97692 80434 97748 80444
rect 97804 80612 97860 80622
rect 97804 80498 97860 80556
rect 97804 80446 97806 80498
rect 97858 80446 97860 80498
rect 97804 80434 97860 80446
rect 97580 79604 97636 79614
rect 97580 79510 97636 79548
rect 97804 78930 97860 78942
rect 97804 78878 97806 78930
rect 97858 78878 97860 78930
rect 97804 78596 97860 78878
rect 97804 78530 97860 78540
rect 97804 75570 97860 75582
rect 97804 75518 97806 75570
rect 97858 75518 97860 75570
rect 97804 74228 97860 75518
rect 97804 74134 97860 74172
rect 98252 75124 98308 75134
rect 97580 73332 97636 73342
rect 97580 73238 97636 73276
rect 97692 72548 97748 72558
rect 97692 70196 97748 72492
rect 97692 69410 97748 70140
rect 97692 69358 97694 69410
rect 97746 69358 97748 69410
rect 97692 69346 97748 69358
rect 98028 67844 98084 67854
rect 97580 66946 97636 66958
rect 97580 66894 97582 66946
rect 97634 66894 97636 66946
rect 97580 66836 97636 66894
rect 97580 66770 97636 66780
rect 97468 66434 97524 66444
rect 97580 66386 97636 66398
rect 98028 66388 98084 67788
rect 97580 66334 97582 66386
rect 97634 66334 97636 66386
rect 96012 65490 96180 65492
rect 96012 65438 96126 65490
rect 96178 65438 96180 65490
rect 96012 65436 96180 65438
rect 96012 63922 96068 65436
rect 96124 65426 96180 65436
rect 96348 65604 96404 65614
rect 96348 65268 96404 65548
rect 97580 65604 97636 66334
rect 97580 65538 97636 65548
rect 97692 66386 98084 66388
rect 97692 66334 98030 66386
rect 98082 66334 98084 66386
rect 97692 66332 98084 66334
rect 96124 65212 96404 65268
rect 96124 64034 96180 65212
rect 96636 65100 96900 65110
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96636 65034 96900 65044
rect 97692 64818 97748 66332
rect 98028 66322 98084 66332
rect 97692 64766 97694 64818
rect 97746 64766 97748 64818
rect 97132 64708 97188 64718
rect 97132 64614 97188 64652
rect 97692 64708 97748 64766
rect 97692 64642 97748 64652
rect 96348 64594 96404 64606
rect 96348 64542 96350 64594
rect 96402 64542 96404 64594
rect 96348 64148 96404 64542
rect 96348 64082 96404 64092
rect 96124 63982 96126 64034
rect 96178 63982 96180 64034
rect 96124 63970 96180 63982
rect 96012 63870 96014 63922
rect 96066 63870 96068 63922
rect 96012 63252 96068 63870
rect 96636 63532 96900 63542
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96636 63466 96900 63476
rect 96124 63252 96180 63262
rect 96012 63250 96180 63252
rect 96012 63198 96126 63250
rect 96178 63198 96180 63250
rect 96012 63196 96180 63198
rect 96124 63186 96180 63196
rect 96460 63140 96516 63150
rect 95788 60734 95790 60786
rect 95842 60734 95844 60786
rect 95788 60722 95844 60734
rect 96348 62356 96404 62366
rect 96348 60116 96404 62300
rect 96460 62242 96516 63084
rect 96460 62190 96462 62242
rect 96514 62190 96516 62242
rect 96460 62178 96516 62190
rect 97020 62916 97076 62926
rect 96636 61964 96900 61974
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96636 61898 96900 61908
rect 96796 61684 96852 61694
rect 97020 61684 97076 62860
rect 96796 61682 97076 61684
rect 96796 61630 96798 61682
rect 96850 61630 97076 61682
rect 96796 61628 97076 61630
rect 97244 62692 97300 62702
rect 96796 61618 96852 61628
rect 96636 60396 96900 60406
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96636 60330 96900 60340
rect 96460 60116 96516 60126
rect 96348 60114 97188 60116
rect 96348 60062 96462 60114
rect 96514 60062 97188 60114
rect 96348 60060 97188 60062
rect 96460 60050 96516 60060
rect 97020 59890 97076 59902
rect 97020 59838 97022 59890
rect 97074 59838 97076 59890
rect 97020 59668 97076 59838
rect 97132 59890 97188 60060
rect 97132 59838 97134 59890
rect 97186 59838 97188 59890
rect 97132 59826 97188 59838
rect 97244 59668 97300 62636
rect 98140 60788 98196 60798
rect 97692 60004 97748 60014
rect 97692 59910 97748 59948
rect 97356 59892 97412 59902
rect 97356 59798 97412 59836
rect 98028 59892 98084 59902
rect 98028 59798 98084 59836
rect 97916 59780 97972 59790
rect 97020 59612 97300 59668
rect 97580 59778 97972 59780
rect 97580 59726 97918 59778
rect 97970 59726 97972 59778
rect 97580 59724 97972 59726
rect 97132 59442 97188 59612
rect 97132 59390 97134 59442
rect 97186 59390 97188 59442
rect 97132 59378 97188 59390
rect 95564 59332 95620 59342
rect 95564 58436 95620 59276
rect 95788 59330 95844 59342
rect 95788 59278 95790 59330
rect 95842 59278 95844 59330
rect 95676 58436 95732 58446
rect 95564 58434 95732 58436
rect 95564 58382 95678 58434
rect 95730 58382 95732 58434
rect 95564 58380 95732 58382
rect 95676 58370 95732 58380
rect 95564 58210 95620 58222
rect 95564 58158 95566 58210
rect 95618 58158 95620 58210
rect 95564 56644 95620 58158
rect 95788 57652 95844 59278
rect 95900 59218 95956 59230
rect 95900 59166 95902 59218
rect 95954 59166 95956 59218
rect 95900 59108 95956 59166
rect 96348 59108 96404 59118
rect 95900 59106 96516 59108
rect 95900 59054 96350 59106
rect 96402 59054 96516 59106
rect 95900 59052 96516 59054
rect 96348 59042 96404 59052
rect 96460 58322 96516 59052
rect 96636 58828 96900 58838
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96636 58762 96900 58772
rect 96460 58270 96462 58322
rect 96514 58270 96516 58322
rect 96124 58210 96180 58222
rect 96124 58158 96126 58210
rect 96178 58158 96180 58210
rect 96124 57876 96180 58158
rect 96124 57810 96180 57820
rect 96348 58210 96404 58222
rect 96348 58158 96350 58210
rect 96402 58158 96404 58210
rect 96348 57764 96404 58158
rect 96460 58100 96516 58270
rect 97580 58324 97636 59724
rect 97916 59714 97972 59724
rect 96460 58034 96516 58044
rect 96908 58210 96964 58222
rect 96908 58158 96910 58210
rect 96962 58158 96964 58210
rect 96908 58100 96964 58158
rect 97356 58210 97412 58222
rect 97356 58158 97358 58210
rect 97410 58158 97412 58210
rect 97356 58100 97412 58158
rect 96908 58034 96964 58044
rect 97244 58044 97356 58100
rect 96348 57708 97188 57764
rect 95788 57596 96516 57652
rect 96460 57538 96516 57596
rect 96460 57486 96462 57538
rect 96514 57486 96516 57538
rect 96460 57474 96516 57486
rect 96636 57260 96900 57270
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96636 57194 96900 57204
rect 97132 56978 97188 57708
rect 97244 57762 97300 58044
rect 97356 58034 97412 58044
rect 97580 57874 97636 58268
rect 97580 57822 97582 57874
rect 97634 57822 97636 57874
rect 97580 57810 97636 57822
rect 97244 57710 97246 57762
rect 97298 57710 97300 57762
rect 97244 57698 97300 57710
rect 97356 57762 97412 57774
rect 97356 57710 97358 57762
rect 97410 57710 97412 57762
rect 97356 57652 97412 57710
rect 97356 57596 97524 57652
rect 97468 57204 97524 57596
rect 97132 56926 97134 56978
rect 97186 56926 97188 56978
rect 97132 56914 97188 56926
rect 97244 57148 97524 57204
rect 97916 57538 97972 57550
rect 97916 57486 97918 57538
rect 97970 57486 97972 57538
rect 97244 56644 97300 57148
rect 95564 56578 95620 56588
rect 96460 56588 97300 56644
rect 97580 56644 97636 56654
rect 97916 56644 97972 57486
rect 97580 56642 97972 56644
rect 97580 56590 97582 56642
rect 97634 56590 97972 56642
rect 97580 56588 97972 56590
rect 96236 55970 96292 55982
rect 96236 55918 96238 55970
rect 96290 55918 96292 55970
rect 96236 55860 96292 55918
rect 96236 55794 96292 55804
rect 94668 54738 94836 54740
rect 94668 54686 94670 54738
rect 94722 54686 94836 54738
rect 94668 54684 94836 54686
rect 95228 55412 95508 55468
rect 94668 54674 94724 54684
rect 93548 54574 93550 54626
rect 93602 54574 93604 54626
rect 92876 53890 92932 53900
rect 93100 53956 93156 53966
rect 93100 53842 93156 53900
rect 93100 53790 93102 53842
rect 93154 53790 93156 53842
rect 93100 53778 93156 53790
rect 93548 53844 93604 54574
rect 93660 54628 93716 54638
rect 93660 54068 93716 54572
rect 94444 54626 94500 54638
rect 94444 54574 94446 54626
rect 94498 54574 94500 54626
rect 93660 54002 93716 54012
rect 94332 54514 94388 54526
rect 94332 54462 94334 54514
rect 94386 54462 94388 54514
rect 93660 53844 93716 53854
rect 94108 53844 94164 53854
rect 94332 53844 94388 54462
rect 94444 54292 94500 54574
rect 94444 54226 94500 54236
rect 95004 54402 95060 54414
rect 95004 54350 95006 54402
rect 95058 54350 95060 54402
rect 95004 54292 95060 54350
rect 95004 54226 95060 54236
rect 93548 53842 94388 53844
rect 93548 53790 93662 53842
rect 93714 53790 94110 53842
rect 94162 53790 94388 53842
rect 93548 53788 94388 53790
rect 94780 53842 94836 53854
rect 94780 53790 94782 53842
rect 94834 53790 94836 53842
rect 93660 53778 93716 53788
rect 94108 53778 94164 53788
rect 94780 53732 94836 53790
rect 94780 53666 94836 53676
rect 94108 53620 94164 53630
rect 92652 53004 92820 53060
rect 92652 52836 92708 52846
rect 92540 52834 92708 52836
rect 92540 52782 92654 52834
rect 92706 52782 92708 52834
rect 92540 52780 92708 52782
rect 92652 52770 92708 52780
rect 92428 52164 92484 52174
rect 92428 52162 92596 52164
rect 92428 52110 92430 52162
rect 92482 52110 92596 52162
rect 92428 52108 92596 52110
rect 92428 52098 92484 52108
rect 91980 51326 91982 51378
rect 92034 51326 92036 51378
rect 91868 50708 91924 50718
rect 91868 50484 91924 50652
rect 91868 50390 91924 50428
rect 91756 50318 91758 50370
rect 91810 50318 91812 50370
rect 91308 50204 91588 50260
rect 91196 49698 91252 49980
rect 91196 49646 91198 49698
rect 91250 49646 91252 49698
rect 91196 49634 91252 49646
rect 90972 47506 91028 47516
rect 90076 45838 90078 45890
rect 90130 45838 90132 45890
rect 90076 45826 90132 45838
rect 90412 46284 90692 46340
rect 91420 46900 91476 46910
rect 89852 45726 89854 45778
rect 89906 45726 89908 45778
rect 89852 45714 89908 45726
rect 89628 45602 89684 45612
rect 90076 44100 90132 44110
rect 89740 43428 89796 43438
rect 89740 43426 89908 43428
rect 89740 43374 89742 43426
rect 89794 43374 89908 43426
rect 89740 43372 89908 43374
rect 89740 43362 89796 43372
rect 89740 42756 89796 42766
rect 89740 42662 89796 42700
rect 89292 42532 89348 42542
rect 89292 41970 89348 42476
rect 89292 41918 89294 41970
rect 89346 41918 89348 41970
rect 89292 41906 89348 41918
rect 89404 42530 89460 42542
rect 89404 42478 89406 42530
rect 89458 42478 89460 42530
rect 89292 40628 89348 40638
rect 89292 40534 89348 40572
rect 89404 40404 89460 42478
rect 89740 41412 89796 41422
rect 89628 41188 89684 41198
rect 89628 41094 89684 41132
rect 89516 40404 89572 40414
rect 89404 40402 89572 40404
rect 89404 40350 89518 40402
rect 89570 40350 89572 40402
rect 89404 40348 89572 40350
rect 89516 40338 89572 40348
rect 89740 39844 89796 41356
rect 89852 41300 89908 43372
rect 90076 43426 90132 44044
rect 90412 43708 90468 46284
rect 90860 46004 90916 46014
rect 90524 45892 90580 45902
rect 90524 45798 90580 45836
rect 90860 45890 90916 45948
rect 91308 46004 91364 46014
rect 91308 45910 91364 45948
rect 90860 45838 90862 45890
rect 90914 45838 90916 45890
rect 90860 45826 90916 45838
rect 91196 45892 91252 45902
rect 90748 45780 90804 45790
rect 90748 45686 90804 45724
rect 91196 44210 91252 45836
rect 91420 45106 91476 46844
rect 91420 45054 91422 45106
rect 91474 45054 91476 45106
rect 91196 44158 91198 44210
rect 91250 44158 91252 44210
rect 91196 44146 91252 44158
rect 91308 44322 91364 44334
rect 91308 44270 91310 44322
rect 91362 44270 91364 44322
rect 90636 44100 90692 44110
rect 90636 44006 90692 44044
rect 91308 44100 91364 44270
rect 90076 43374 90078 43426
rect 90130 43374 90132 43426
rect 90076 42868 90132 43374
rect 90076 42802 90132 42812
rect 90188 43652 90468 43708
rect 89964 42642 90020 42654
rect 89964 42590 89966 42642
rect 90018 42590 90020 42642
rect 89964 42196 90020 42590
rect 89964 42130 90020 42140
rect 89852 41234 89908 41244
rect 90188 41076 90244 43652
rect 90524 42642 90580 42654
rect 90524 42590 90526 42642
rect 90578 42590 90580 42642
rect 90300 41412 90356 41422
rect 90524 41412 90580 42590
rect 90524 41356 91140 41412
rect 90300 41318 90356 41356
rect 90412 41300 90468 41310
rect 90468 41244 90692 41300
rect 90412 41234 90468 41244
rect 90636 41186 90692 41244
rect 90636 41134 90638 41186
rect 90690 41134 90692 41186
rect 90188 41020 90468 41076
rect 89404 39788 89796 39844
rect 89404 38834 89460 39788
rect 90076 39508 90132 39518
rect 89628 39506 90132 39508
rect 89628 39454 90078 39506
rect 90130 39454 90132 39506
rect 89628 39452 90132 39454
rect 89628 39058 89684 39452
rect 90076 39442 90132 39452
rect 89628 39006 89630 39058
rect 89682 39006 89684 39058
rect 89628 38994 89684 39006
rect 89404 38782 89406 38834
rect 89458 38782 89460 38834
rect 89404 38770 89460 38782
rect 90188 38948 90244 38958
rect 90188 38834 90244 38892
rect 90188 38782 90190 38834
rect 90242 38782 90244 38834
rect 89180 38220 89348 38276
rect 89180 38050 89236 38062
rect 89180 37998 89182 38050
rect 89234 37998 89236 38050
rect 89180 36708 89236 37998
rect 89292 37156 89348 38220
rect 89516 38052 89572 38062
rect 89404 37826 89460 37838
rect 89404 37774 89406 37826
rect 89458 37774 89460 37826
rect 89404 37380 89460 37774
rect 89404 37314 89460 37324
rect 89292 37024 89348 37100
rect 89180 36652 89460 36708
rect 88732 36530 88788 36540
rect 89404 35922 89460 36652
rect 89516 36596 89572 37996
rect 89852 37828 89908 37838
rect 90188 37828 90244 38782
rect 89852 37826 90244 37828
rect 89852 37774 89854 37826
rect 89906 37774 90244 37826
rect 89852 37772 90244 37774
rect 89516 36594 89796 36596
rect 89516 36542 89518 36594
rect 89570 36542 89796 36594
rect 89516 36540 89796 36542
rect 89516 36530 89572 36540
rect 89404 35870 89406 35922
rect 89458 35870 89460 35922
rect 89404 35858 89460 35870
rect 88508 35812 88564 35822
rect 88508 35028 88564 35756
rect 89740 35698 89796 36540
rect 89740 35646 89742 35698
rect 89794 35646 89796 35698
rect 89740 35634 89796 35646
rect 89852 35476 89908 37772
rect 90300 37156 90356 37166
rect 89964 35812 90020 35822
rect 89964 35718 90020 35756
rect 90300 35810 90356 37100
rect 90300 35758 90302 35810
rect 90354 35758 90356 35810
rect 89628 35420 89908 35476
rect 88620 35028 88676 35038
rect 88508 35026 88676 35028
rect 88508 34974 88622 35026
rect 88674 34974 88676 35026
rect 88508 34972 88676 34974
rect 88620 34962 88676 34972
rect 89516 34916 89572 34926
rect 88396 34066 88452 34076
rect 88620 34692 88676 34702
rect 88620 33458 88676 34636
rect 88620 33406 88622 33458
rect 88674 33406 88676 33458
rect 88508 32788 88564 32798
rect 88620 32788 88676 33406
rect 88172 32722 88228 32732
rect 88284 32786 88676 32788
rect 88284 32734 88510 32786
rect 88562 32734 88676 32786
rect 88284 32732 88676 32734
rect 89180 34132 89236 34142
rect 89180 32786 89236 34076
rect 89404 34132 89460 34142
rect 89404 34038 89460 34076
rect 89516 33684 89572 34860
rect 89516 33458 89572 33628
rect 89516 33406 89518 33458
rect 89570 33406 89572 33458
rect 89516 33394 89572 33406
rect 89180 32734 89182 32786
rect 89234 32734 89236 32786
rect 87388 32676 87444 32686
rect 87388 32582 87444 32620
rect 87836 32674 87892 32686
rect 87836 32622 87838 32674
rect 87890 32622 87892 32674
rect 87836 32564 87892 32622
rect 88284 32564 88340 32732
rect 88508 32722 88564 32732
rect 89180 32722 89236 32734
rect 87836 32508 88340 32564
rect 86940 31838 86942 31890
rect 86994 31838 86996 31890
rect 86940 31826 86996 31838
rect 87052 32338 87108 32350
rect 87052 32286 87054 32338
rect 87106 32286 87108 32338
rect 86044 30884 86100 30894
rect 86044 30790 86100 30828
rect 87052 30884 87108 32286
rect 89292 31892 89348 31902
rect 89292 31798 89348 31836
rect 87052 30818 87108 30828
rect 85428 29372 85652 29428
rect 85372 29296 85428 29372
rect 81676 8372 81956 8428
rect 82460 8372 82628 8428
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 80780 3444 80836 3454
rect 81228 3444 81284 3454
rect 80780 3442 81284 3444
rect 80780 3390 80782 3442
rect 80834 3390 81230 3442
rect 81282 3390 81284 3442
rect 80780 3388 81284 3390
rect 80780 3378 80836 3388
rect 77532 2818 77588 2828
rect 69020 2706 69076 2716
rect 68572 2268 68852 2324
rect 68572 800 68628 2268
rect 81004 800 81060 3388
rect 81228 3378 81284 3388
rect 81564 3332 81620 3342
rect 81676 3332 81732 8372
rect 81564 3330 81732 3332
rect 81564 3278 81566 3330
rect 81618 3278 81732 3330
rect 81564 3276 81732 3278
rect 81564 3266 81620 3276
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 82460 2996 82516 8372
rect 89628 3332 89684 35420
rect 90300 35026 90356 35758
rect 90412 35308 90468 41020
rect 90636 39732 90692 41134
rect 90748 41188 90804 41198
rect 90748 40292 90804 41132
rect 91084 41076 91140 41356
rect 91308 41188 91364 44044
rect 91420 43540 91476 45054
rect 91420 43474 91476 43484
rect 91196 41076 91252 41086
rect 91084 41074 91252 41076
rect 91084 41022 91198 41074
rect 91250 41022 91252 41074
rect 91308 41056 91364 41132
rect 91084 41020 91252 41022
rect 90860 40292 90916 40302
rect 90748 40290 90916 40292
rect 90748 40238 90862 40290
rect 90914 40238 90916 40290
rect 90748 40236 90916 40238
rect 90636 39666 90692 39676
rect 90860 39618 90916 40236
rect 90860 39566 90862 39618
rect 90914 39566 90916 39618
rect 90860 39554 90916 39566
rect 90524 38948 90580 38958
rect 91084 38948 91140 41020
rect 91196 41010 91252 41020
rect 90524 38946 91140 38948
rect 90524 38894 90526 38946
rect 90578 38894 91140 38946
rect 90524 38892 91140 38894
rect 91532 38948 91588 50204
rect 91756 49700 91812 50318
rect 91756 49634 91812 49644
rect 91980 49026 92036 51326
rect 92428 50596 92484 50606
rect 92428 50502 92484 50540
rect 92540 50484 92596 52108
rect 92540 50418 92596 50428
rect 91980 48974 91982 49026
rect 92034 48974 92036 49026
rect 91980 46900 92036 48974
rect 92652 49812 92708 49822
rect 92652 48466 92708 49756
rect 92652 48414 92654 48466
rect 92706 48414 92708 48466
rect 92652 48402 92708 48414
rect 92204 48356 92260 48366
rect 92204 48130 92260 48300
rect 92204 48078 92206 48130
rect 92258 48078 92260 48130
rect 92204 48066 92260 48078
rect 92092 47572 92148 47582
rect 92092 47478 92148 47516
rect 91980 46834 92036 46844
rect 92540 46562 92596 46574
rect 92540 46510 92542 46562
rect 92594 46510 92596 46562
rect 92428 46004 92484 46014
rect 92428 45910 92484 45948
rect 92540 45780 92596 46510
rect 92540 45714 92596 45724
rect 91980 45668 92036 45678
rect 91980 45218 92036 45612
rect 91980 45166 91982 45218
rect 92034 45166 92036 45218
rect 91980 45154 92036 45166
rect 91980 44324 92036 44334
rect 91980 44230 92036 44268
rect 92316 44098 92372 44110
rect 92316 44046 92318 44098
rect 92370 44046 92372 44098
rect 92316 42756 92372 44046
rect 92764 43708 92820 53004
rect 93996 52948 94052 52958
rect 93212 52834 93268 52846
rect 93212 52782 93214 52834
rect 93266 52782 93268 52834
rect 93212 52052 93268 52782
rect 93548 52836 93604 52846
rect 93996 52836 94052 52892
rect 93548 52834 94052 52836
rect 93548 52782 93550 52834
rect 93602 52782 93998 52834
rect 94050 52782 94052 52834
rect 93548 52780 94052 52782
rect 93548 52770 93604 52780
rect 93324 52220 93604 52276
rect 93324 52052 93380 52220
rect 93212 52050 93380 52052
rect 93212 51998 93326 52050
rect 93378 51998 93380 52050
rect 93212 51996 93380 51998
rect 93324 51986 93380 51996
rect 93436 52050 93492 52062
rect 93436 51998 93438 52050
rect 93490 51998 93492 52050
rect 93100 51938 93156 51950
rect 93100 51886 93102 51938
rect 93154 51886 93156 51938
rect 92988 50596 93044 50606
rect 92876 48356 92932 48366
rect 92876 48262 92932 48300
rect 92988 48354 93044 50540
rect 93100 50260 93156 51886
rect 93212 51604 93268 51614
rect 93212 50596 93268 51548
rect 93324 50820 93380 50830
rect 93436 50820 93492 51998
rect 93324 50818 93492 50820
rect 93324 50766 93326 50818
rect 93378 50766 93492 50818
rect 93324 50764 93492 50766
rect 93324 50754 93380 50764
rect 93212 50594 93492 50596
rect 93212 50542 93214 50594
rect 93266 50542 93492 50594
rect 93212 50540 93492 50542
rect 93212 50530 93268 50540
rect 93324 50372 93380 50382
rect 93324 50278 93380 50316
rect 93100 50204 93268 50260
rect 93212 49924 93268 50204
rect 93324 49924 93380 49934
rect 93212 49922 93380 49924
rect 93212 49870 93326 49922
rect 93378 49870 93380 49922
rect 93212 49868 93380 49870
rect 93324 49858 93380 49868
rect 93436 49700 93492 50540
rect 93212 49644 93492 49700
rect 93212 49138 93268 49644
rect 93212 49086 93214 49138
rect 93266 49086 93268 49138
rect 93212 49074 93268 49086
rect 93548 48916 93604 52220
rect 93996 52050 94052 52780
rect 93996 51998 93998 52050
rect 94050 51998 94052 52050
rect 93996 51604 94052 51998
rect 94108 52050 94164 53564
rect 94668 53060 94724 53070
rect 94668 52966 94724 53004
rect 94556 52948 94612 52958
rect 94556 52854 94612 52892
rect 94668 52722 94724 52734
rect 94668 52670 94670 52722
rect 94722 52670 94724 52722
rect 94332 52164 94388 52174
rect 94332 52070 94388 52108
rect 94108 51998 94110 52050
rect 94162 51998 94164 52050
rect 94108 51986 94164 51998
rect 93996 51538 94052 51548
rect 94108 51828 94164 51838
rect 93996 51156 94052 51166
rect 93996 50594 94052 51100
rect 93996 50542 93998 50594
rect 94050 50542 94052 50594
rect 93884 50484 93940 50494
rect 92988 48302 92990 48354
rect 93042 48302 93044 48354
rect 92988 46004 93044 48302
rect 93100 48860 93604 48916
rect 93772 48916 93828 48926
rect 93100 46786 93156 48860
rect 93772 48822 93828 48860
rect 93660 48244 93716 48254
rect 93660 48150 93716 48188
rect 93436 48132 93492 48142
rect 93212 47348 93268 47358
rect 93212 47254 93268 47292
rect 93324 47236 93380 47246
rect 93212 46900 93268 46910
rect 93324 46900 93380 47180
rect 93212 46898 93380 46900
rect 93212 46846 93214 46898
rect 93266 46846 93380 46898
rect 93212 46844 93380 46846
rect 93436 46898 93492 48076
rect 93548 47460 93604 47470
rect 93548 47346 93604 47404
rect 93548 47294 93550 47346
rect 93602 47294 93604 47346
rect 93548 47282 93604 47294
rect 93660 47348 93716 47358
rect 93436 46846 93438 46898
rect 93490 46846 93492 46898
rect 93212 46834 93268 46844
rect 93436 46834 93492 46846
rect 93100 46734 93102 46786
rect 93154 46734 93156 46786
rect 93100 46452 93156 46734
rect 93100 46386 93156 46396
rect 93660 46564 93716 47292
rect 93884 47012 93940 50428
rect 93996 50260 94052 50542
rect 94108 50482 94164 51772
rect 94668 51604 94724 52670
rect 94892 52724 94948 52734
rect 94780 52276 94836 52286
rect 94892 52276 94948 52668
rect 94780 52274 94948 52276
rect 94780 52222 94782 52274
rect 94834 52222 94948 52274
rect 94780 52220 94948 52222
rect 94780 52210 94836 52220
rect 94668 51538 94724 51548
rect 95004 51492 95060 51502
rect 95004 50596 95060 51436
rect 94108 50430 94110 50482
rect 94162 50430 94164 50482
rect 94108 50418 94164 50430
rect 94220 50594 95060 50596
rect 94220 50542 95006 50594
rect 95058 50542 95060 50594
rect 94220 50540 95060 50542
rect 94108 50260 94164 50270
rect 93996 50204 94108 50260
rect 94108 50194 94164 50204
rect 94108 49812 94164 49822
rect 94220 49812 94276 50540
rect 95004 50530 95060 50540
rect 94332 50372 94388 50382
rect 94332 50278 94388 50316
rect 94892 50260 94948 50270
rect 94780 49922 94836 49934
rect 94780 49870 94782 49922
rect 94834 49870 94836 49922
rect 94108 49810 94276 49812
rect 94108 49758 94110 49810
rect 94162 49758 94276 49810
rect 94108 49756 94276 49758
rect 94108 49746 94164 49756
rect 94108 48914 94164 48926
rect 94108 48862 94110 48914
rect 94162 48862 94164 48914
rect 94108 47348 94164 48862
rect 94220 48244 94276 49756
rect 94220 48178 94276 48188
rect 94556 49810 94612 49822
rect 94556 49758 94558 49810
rect 94610 49758 94612 49810
rect 94332 48132 94388 48142
rect 94332 48038 94388 48076
rect 94444 48020 94500 48030
rect 94108 47282 94164 47292
rect 94332 47346 94388 47358
rect 94332 47294 94334 47346
rect 94386 47294 94388 47346
rect 93996 47234 94052 47246
rect 93996 47182 93998 47234
rect 94050 47182 94052 47234
rect 93996 47124 94052 47182
rect 93996 47058 94052 47068
rect 94220 47234 94276 47246
rect 94220 47182 94222 47234
rect 94274 47182 94276 47234
rect 94220 47124 94276 47182
rect 93884 46946 93940 46956
rect 93772 46900 93828 46910
rect 93772 46806 93828 46844
rect 92988 45938 93044 45948
rect 93324 45892 93380 45902
rect 93100 45668 93156 45678
rect 93100 44434 93156 45612
rect 93100 44382 93102 44434
rect 93154 44382 93156 44434
rect 92764 43652 92932 43708
rect 92316 42690 92372 42700
rect 92652 43540 92708 43550
rect 92428 42532 92484 42542
rect 92428 42438 92484 42476
rect 92652 42084 92708 43484
rect 92652 41860 92708 42028
rect 92652 41794 92708 41804
rect 92428 41076 92484 41086
rect 92428 40982 92484 41020
rect 92092 40964 92148 40974
rect 90524 38882 90580 38892
rect 90860 37938 90916 38892
rect 91532 38882 91588 38892
rect 91868 40962 92148 40964
rect 91868 40910 92094 40962
rect 92146 40910 92148 40962
rect 91868 40908 92148 40910
rect 91868 38946 91924 40908
rect 92092 40898 92148 40908
rect 91868 38894 91870 38946
rect 91922 38894 91924 38946
rect 91868 38882 91924 38894
rect 91196 38836 91252 38846
rect 91196 38742 91252 38780
rect 90860 37886 90862 37938
rect 90914 37886 90916 37938
rect 90412 35252 90804 35308
rect 90300 34974 90302 35026
rect 90354 34974 90356 35026
rect 90300 34962 90356 34974
rect 89852 34690 89908 34702
rect 89852 34638 89854 34690
rect 89906 34638 89908 34690
rect 89852 34356 89908 34638
rect 89852 34290 89908 34300
rect 90076 34018 90132 34030
rect 90076 33966 90078 34018
rect 90130 33966 90132 34018
rect 89852 32338 89908 32350
rect 89852 32286 89854 32338
rect 89906 32286 89908 32338
rect 89852 31778 89908 32286
rect 89852 31726 89854 31778
rect 89906 31726 89908 31778
rect 89852 31714 89908 31726
rect 90076 31666 90132 33966
rect 90748 34020 90804 35252
rect 90860 34802 90916 37886
rect 90972 38050 91028 38062
rect 90972 37998 90974 38050
rect 91026 37998 91028 38050
rect 90972 37828 91028 37998
rect 91644 38052 91700 38062
rect 91644 37958 91700 37996
rect 90972 36596 91028 37772
rect 91980 37826 92036 37838
rect 91980 37774 91982 37826
rect 92034 37774 92036 37826
rect 91420 37380 91476 37390
rect 91420 37286 91476 37324
rect 91980 37380 92036 37774
rect 91980 37314 92036 37324
rect 92764 37378 92820 37390
rect 92764 37326 92766 37378
rect 92818 37326 92820 37378
rect 92204 37266 92260 37278
rect 92204 37214 92206 37266
rect 92258 37214 92260 37266
rect 90972 36530 91028 36540
rect 91644 37044 91700 37054
rect 91644 36594 91700 36988
rect 91644 36542 91646 36594
rect 91698 36542 91700 36594
rect 91644 36530 91700 36542
rect 92204 36484 92260 37214
rect 92764 37044 92820 37326
rect 92764 36978 92820 36988
rect 92428 36484 92484 36494
rect 92204 36482 92484 36484
rect 92204 36430 92430 36482
rect 92482 36430 92484 36482
rect 92204 36428 92484 36430
rect 90860 34750 90862 34802
rect 90914 34750 90916 34802
rect 90860 34738 90916 34750
rect 90972 34914 91028 34926
rect 90972 34862 90974 34914
rect 91026 34862 91028 34914
rect 90972 34468 91028 34862
rect 91644 34916 91700 34926
rect 91644 34822 91700 34860
rect 90972 34402 91028 34412
rect 91980 34690 92036 34702
rect 91980 34638 91982 34690
rect 92034 34638 92036 34690
rect 91980 34244 92036 34638
rect 91980 34178 92036 34188
rect 92428 34132 92484 36428
rect 92876 35252 92932 43652
rect 92988 42196 93044 42206
rect 92988 38612 93044 42140
rect 93100 38836 93156 44382
rect 93324 44546 93380 45836
rect 93548 45668 93604 45678
rect 93660 45668 93716 46508
rect 94108 46004 94164 46014
rect 94220 46004 94276 47068
rect 94332 47012 94388 47294
rect 94332 46946 94388 46956
rect 94332 46562 94388 46574
rect 94332 46510 94334 46562
rect 94386 46510 94388 46562
rect 94332 46114 94388 46510
rect 94332 46062 94334 46114
rect 94386 46062 94388 46114
rect 94332 46050 94388 46062
rect 94108 46002 94276 46004
rect 94108 45950 94110 46002
rect 94162 45950 94276 46002
rect 94108 45948 94276 45950
rect 94108 45938 94164 45948
rect 93548 45666 93828 45668
rect 93548 45614 93550 45666
rect 93602 45614 93828 45666
rect 93548 45612 93828 45614
rect 93548 45602 93604 45612
rect 93324 44494 93326 44546
rect 93378 44494 93380 44546
rect 93212 42756 93268 42766
rect 93212 42662 93268 42700
rect 93212 41300 93268 41310
rect 93324 41300 93380 44494
rect 93548 44324 93604 44334
rect 93548 43708 93604 44268
rect 93548 43652 93716 43708
rect 93212 41298 93380 41300
rect 93212 41246 93214 41298
rect 93266 41246 93380 41298
rect 93212 41244 93380 41246
rect 93548 42530 93604 42542
rect 93548 42478 93550 42530
rect 93602 42478 93604 42530
rect 93548 41300 93604 42478
rect 93212 41234 93268 41244
rect 93548 41234 93604 41244
rect 93660 40516 93716 43652
rect 93660 40450 93716 40460
rect 93324 39732 93380 39742
rect 93772 39732 93828 45612
rect 94444 45444 94500 47964
rect 94556 47236 94612 49758
rect 94780 49700 94836 49870
rect 94892 49924 94948 50204
rect 94892 49792 94948 49868
rect 94780 49634 94836 49644
rect 94892 49138 94948 49150
rect 94892 49086 94894 49138
rect 94946 49086 94948 49138
rect 94780 48244 94836 48254
rect 94780 47572 94836 48188
rect 94892 47796 94948 49086
rect 95228 48916 95284 55412
rect 96460 55410 96516 56588
rect 97244 55972 97300 55982
rect 97244 55878 97300 55916
rect 97020 55860 97076 55870
rect 96636 55692 96900 55702
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96636 55626 96900 55636
rect 96460 55358 96462 55410
rect 96514 55358 96516 55410
rect 96460 55346 96516 55358
rect 96908 55412 96964 55422
rect 97020 55412 97076 55804
rect 97580 55860 97636 56588
rect 97580 55794 97636 55804
rect 97804 55972 97860 55982
rect 96908 55410 97076 55412
rect 96908 55358 96910 55410
rect 96962 55358 97076 55410
rect 96908 55356 97076 55358
rect 96908 55346 96964 55356
rect 95564 54292 95620 54302
rect 95452 53058 95508 53070
rect 95452 53006 95454 53058
rect 95506 53006 95508 53058
rect 95340 52946 95396 52958
rect 95340 52894 95342 52946
rect 95394 52894 95396 52946
rect 95340 52164 95396 52894
rect 95340 52098 95396 52108
rect 95452 50148 95508 53006
rect 95452 50082 95508 50092
rect 95564 50034 95620 54236
rect 96636 54124 96900 54134
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96636 54058 96900 54068
rect 97692 53732 97748 53742
rect 96908 53618 96964 53630
rect 96908 53566 96910 53618
rect 96962 53566 96964 53618
rect 95676 53172 95732 53182
rect 95676 53078 95732 53116
rect 96908 53172 96964 53566
rect 96908 53106 96964 53116
rect 96236 53058 96292 53070
rect 96236 53006 96238 53058
rect 96290 53006 96292 53058
rect 96124 52948 96180 52958
rect 96124 52612 96180 52892
rect 95564 49982 95566 50034
rect 95618 49982 95620 50034
rect 95452 49924 95508 49934
rect 95452 49830 95508 49868
rect 95228 48850 95284 48860
rect 95340 49700 95396 49710
rect 94892 47730 94948 47740
rect 94556 47170 94612 47180
rect 94668 47570 95172 47572
rect 94668 47518 94782 47570
rect 94834 47518 95172 47570
rect 94668 47516 95172 47518
rect 94668 46002 94724 47516
rect 94780 47506 94836 47516
rect 95116 46898 95172 47516
rect 95228 47348 95284 47358
rect 95228 47254 95284 47292
rect 95116 46846 95118 46898
rect 95170 46846 95172 46898
rect 95116 46834 95172 46846
rect 94780 46562 94836 46574
rect 94780 46510 94782 46562
rect 94834 46510 94836 46562
rect 94780 46450 94836 46510
rect 94780 46398 94782 46450
rect 94834 46398 94836 46450
rect 94780 46386 94836 46398
rect 95116 46452 95172 46462
rect 94668 45950 94670 46002
rect 94722 45950 94724 46002
rect 94668 45938 94724 45950
rect 95116 46002 95172 46396
rect 95340 46114 95396 49644
rect 95564 47460 95620 49982
rect 95676 50482 95732 50494
rect 95676 50430 95678 50482
rect 95730 50430 95732 50482
rect 95676 50036 95732 50430
rect 96124 50260 96180 52556
rect 96236 51940 96292 53006
rect 96236 51874 96292 51884
rect 96460 52948 96516 52958
rect 97580 52948 97636 52958
rect 96460 52946 97076 52948
rect 96460 52894 96462 52946
rect 96514 52894 97076 52946
rect 96460 52892 97076 52894
rect 96236 51492 96292 51502
rect 96236 51398 96292 51436
rect 96348 50372 96404 50382
rect 96124 50204 96292 50260
rect 95676 49970 95732 49980
rect 96124 50036 96180 50046
rect 96124 49942 96180 49980
rect 95788 49924 95844 49934
rect 95788 49830 95844 49868
rect 95564 46900 95620 47404
rect 95564 46834 95620 46844
rect 95676 49812 95732 49822
rect 95676 46898 95732 49756
rect 96236 48356 96292 50204
rect 96348 50034 96404 50316
rect 96348 49982 96350 50034
rect 96402 49982 96404 50034
rect 96348 49970 96404 49982
rect 96460 49922 96516 52892
rect 96636 52556 96900 52566
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96636 52490 96900 52500
rect 97020 52276 97076 52892
rect 97580 52854 97636 52892
rect 97132 52836 97188 52846
rect 97132 52742 97188 52780
rect 97020 52220 97412 52276
rect 96908 52052 96964 52062
rect 96908 52050 97188 52052
rect 96908 51998 96910 52050
rect 96962 51998 97188 52050
rect 96908 51996 97188 51998
rect 96908 51986 96964 51996
rect 97132 51602 97188 51996
rect 97132 51550 97134 51602
rect 97186 51550 97188 51602
rect 97132 51538 97188 51550
rect 97356 51602 97412 52220
rect 97692 52162 97748 53676
rect 97804 53396 97860 55916
rect 98028 54402 98084 54414
rect 98028 54350 98030 54402
rect 98082 54350 98084 54402
rect 98028 53732 98084 54350
rect 97804 53340 97972 53396
rect 97692 52110 97694 52162
rect 97746 52110 97748 52162
rect 97356 51550 97358 51602
rect 97410 51550 97412 51602
rect 97356 51538 97412 51550
rect 97468 51604 97524 51614
rect 97468 51490 97524 51548
rect 97468 51438 97470 51490
rect 97522 51438 97524 51490
rect 97468 51426 97524 51438
rect 97692 51492 97748 52110
rect 96636 50988 96900 50998
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96636 50922 96900 50932
rect 97468 50148 97524 50158
rect 96460 49870 96462 49922
rect 96514 49870 96516 49922
rect 96460 49858 96516 49870
rect 97356 49924 97412 49934
rect 97356 49830 97412 49868
rect 97468 49924 97524 50092
rect 97468 49922 97636 49924
rect 97468 49870 97470 49922
rect 97522 49870 97636 49922
rect 97468 49868 97636 49870
rect 97468 49858 97524 49868
rect 97132 49810 97188 49822
rect 97132 49758 97134 49810
rect 97186 49758 97188 49810
rect 96636 49420 96900 49430
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96636 49354 96900 49364
rect 97020 49140 97076 49150
rect 97132 49140 97188 49758
rect 97020 49138 97188 49140
rect 97020 49086 97022 49138
rect 97074 49086 97188 49138
rect 97020 49084 97188 49086
rect 97020 49074 97076 49084
rect 97356 48356 97412 48366
rect 96124 48300 96236 48356
rect 96124 47458 96180 48300
rect 96236 48290 96292 48300
rect 96460 48354 97412 48356
rect 96460 48302 97358 48354
rect 97410 48302 97412 48354
rect 96460 48300 97412 48302
rect 96460 48130 96516 48300
rect 97356 48290 97412 48300
rect 97468 48356 97524 48366
rect 97468 48262 97524 48300
rect 96460 48078 96462 48130
rect 96514 48078 96516 48130
rect 96460 48066 96516 48078
rect 97244 48132 97300 48142
rect 96636 47852 96900 47862
rect 96124 47406 96126 47458
rect 96178 47406 96180 47458
rect 96124 47124 96180 47406
rect 96236 47796 96292 47806
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96636 47786 96900 47796
rect 96236 47346 96292 47740
rect 97244 47570 97300 48076
rect 97244 47518 97246 47570
rect 97298 47518 97300 47570
rect 97244 47506 97300 47518
rect 97356 48018 97412 48030
rect 97356 47966 97358 48018
rect 97410 47966 97412 48018
rect 96460 47460 96516 47470
rect 96460 47366 96516 47404
rect 96236 47294 96238 47346
rect 96290 47294 96292 47346
rect 96236 47282 96292 47294
rect 96796 47234 96852 47246
rect 96796 47182 96798 47234
rect 96850 47182 96852 47234
rect 96796 47124 96852 47182
rect 96124 47068 96628 47124
rect 95676 46846 95678 46898
rect 95730 46846 95732 46898
rect 95676 46450 95732 46846
rect 96012 46900 96068 46910
rect 96012 46806 96068 46844
rect 96572 46898 96628 47068
rect 96796 47058 96852 47068
rect 96572 46846 96574 46898
rect 96626 46846 96628 46898
rect 96572 46834 96628 46846
rect 95676 46398 95678 46450
rect 95730 46398 95732 46450
rect 95676 46386 95732 46398
rect 97356 46452 97412 47966
rect 97580 47460 97636 49868
rect 97692 49028 97748 51436
rect 97804 51940 97860 51950
rect 97804 50706 97860 51884
rect 97916 51602 97972 53340
rect 98028 53170 98084 53676
rect 98028 53118 98030 53170
rect 98082 53118 98084 53170
rect 98028 53106 98084 53118
rect 97916 51550 97918 51602
rect 97970 51550 97972 51602
rect 97916 51538 97972 51550
rect 97804 50654 97806 50706
rect 97858 50654 97860 50706
rect 97804 50642 97860 50654
rect 97916 49812 97972 49822
rect 97916 49718 97972 49756
rect 97692 49026 97972 49028
rect 97692 48974 97694 49026
rect 97746 48974 97972 49026
rect 97692 48972 97972 48974
rect 97692 48962 97748 48972
rect 97916 48466 97972 48972
rect 97916 48414 97918 48466
rect 97970 48414 97972 48466
rect 97916 48402 97972 48414
rect 97580 47394 97636 47404
rect 97356 46386 97412 46396
rect 96636 46284 96900 46294
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 95340 46062 95342 46114
rect 95394 46062 95396 46114
rect 95340 46050 95396 46062
rect 95116 45950 95118 46002
rect 95170 45950 95172 46002
rect 95116 45938 95172 45950
rect 95564 45666 95620 45678
rect 95564 45614 95566 45666
rect 95618 45614 95620 45666
rect 94444 45388 94948 45444
rect 93996 44546 94052 44558
rect 93996 44494 93998 44546
rect 94050 44494 94052 44546
rect 93996 44434 94052 44494
rect 93996 44382 93998 44434
rect 94050 44382 94052 44434
rect 93996 44370 94052 44382
rect 94892 44434 94948 45388
rect 94892 44382 94894 44434
rect 94946 44382 94948 44434
rect 94892 43708 94948 44382
rect 94892 43652 95060 43708
rect 94332 42868 94388 42878
rect 94332 42774 94388 42812
rect 94556 42868 94612 42878
rect 94332 41860 94388 41870
rect 94332 41766 94388 41804
rect 93324 39730 93828 39732
rect 93324 39678 93326 39730
rect 93378 39678 93828 39730
rect 93324 39676 93828 39678
rect 93324 39666 93380 39676
rect 93772 39620 93828 39676
rect 93996 40516 94052 40526
rect 93884 39620 93940 39630
rect 93772 39618 93940 39620
rect 93772 39566 93886 39618
rect 93938 39566 93940 39618
rect 93772 39564 93940 39566
rect 93884 39554 93940 39564
rect 93100 38770 93156 38780
rect 93996 38722 94052 40460
rect 94220 39396 94276 39406
rect 94220 39394 94388 39396
rect 94220 39342 94222 39394
rect 94274 39342 94388 39394
rect 94220 39340 94388 39342
rect 94220 39330 94276 39340
rect 93996 38670 93998 38722
rect 94050 38670 94052 38722
rect 93996 38658 94052 38670
rect 94220 38836 94276 38846
rect 93884 38612 93940 38622
rect 92988 38556 93380 38612
rect 93324 38162 93380 38556
rect 93324 38110 93326 38162
rect 93378 38110 93380 38162
rect 93324 38098 93380 38110
rect 93772 37938 93828 37950
rect 93772 37886 93774 37938
rect 93826 37886 93828 37938
rect 93100 37380 93156 37390
rect 93100 37286 93156 37324
rect 93772 36708 93828 37886
rect 93884 37490 93940 38556
rect 94108 37940 94164 37950
rect 94108 37846 94164 37884
rect 93884 37438 93886 37490
rect 93938 37438 93940 37490
rect 93884 37426 93940 37438
rect 94220 37490 94276 38780
rect 94332 38612 94388 39340
rect 94332 38546 94388 38556
rect 94556 39058 94612 42812
rect 94892 42866 94948 42878
rect 94892 42814 94894 42866
rect 94946 42814 94948 42866
rect 94892 41748 94948 42814
rect 95004 42532 95060 43652
rect 95564 43652 95620 45614
rect 95900 45668 95956 45678
rect 95900 45666 96068 45668
rect 95900 45614 95902 45666
rect 95954 45614 96068 45666
rect 95900 45612 96068 45614
rect 95900 45602 95956 45612
rect 95788 45106 95844 45118
rect 95788 45054 95790 45106
rect 95842 45054 95844 45106
rect 95788 44436 95844 45054
rect 95788 44370 95844 44380
rect 96012 44212 96068 45612
rect 96124 45220 96180 45230
rect 96124 45218 97076 45220
rect 96124 45166 96126 45218
rect 96178 45166 97076 45218
rect 96124 45164 97076 45166
rect 96124 45154 96180 45164
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 97020 44434 97076 45164
rect 97020 44382 97022 44434
rect 97074 44382 97076 44434
rect 97020 44370 97076 44382
rect 97692 44322 97748 44334
rect 97692 44270 97694 44322
rect 97746 44270 97748 44322
rect 96012 44156 96292 44212
rect 95900 43876 95956 43886
rect 95564 42868 95620 43596
rect 95564 42802 95620 42812
rect 95788 43764 95844 43774
rect 95004 42466 95060 42476
rect 95340 42532 95396 42542
rect 95340 42082 95396 42476
rect 95340 42030 95342 42082
rect 95394 42030 95396 42082
rect 95340 42018 95396 42030
rect 94892 41682 94948 41692
rect 95228 41972 95284 41982
rect 94892 39732 94948 39742
rect 94892 39638 94948 39676
rect 94556 39006 94558 39058
rect 94610 39006 94612 39058
rect 94556 38052 94612 39006
rect 95228 38834 95284 41916
rect 95676 41860 95732 41870
rect 95788 41860 95844 43708
rect 95900 43708 95956 43820
rect 96236 43764 96292 44156
rect 95900 43652 96068 43708
rect 96236 43698 96292 43708
rect 97020 43764 97076 43774
rect 97020 43652 97188 43708
rect 96012 43092 96068 43652
rect 97132 43650 97188 43652
rect 97132 43598 97134 43650
rect 97186 43598 97188 43650
rect 97132 43586 97188 43598
rect 97692 43652 97748 44270
rect 98140 43708 98196 60732
rect 98252 48020 98308 75068
rect 98252 47954 98308 47964
rect 98140 43652 98308 43708
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96012 43036 96404 43092
rect 96636 43082 96900 43092
rect 95732 41804 95844 41860
rect 96124 42868 96180 42878
rect 95340 41300 95396 41310
rect 95340 41206 95396 41244
rect 95676 40404 95732 41804
rect 96012 41748 96068 41758
rect 95676 40402 95844 40404
rect 95676 40350 95678 40402
rect 95730 40350 95844 40402
rect 95676 40348 95844 40350
rect 95676 40338 95732 40348
rect 95228 38782 95230 38834
rect 95282 38782 95284 38834
rect 95228 38770 95284 38782
rect 95340 39732 95396 39742
rect 94668 38052 94724 38062
rect 94556 38050 94724 38052
rect 94556 37998 94670 38050
rect 94722 37998 94724 38050
rect 94556 37996 94724 37998
rect 94668 37986 94724 37996
rect 94220 37438 94222 37490
rect 94274 37438 94276 37490
rect 94220 37426 94276 37438
rect 95340 37378 95396 39676
rect 95452 38946 95508 38958
rect 95452 38894 95454 38946
rect 95506 38894 95508 38946
rect 95452 38612 95508 38894
rect 95788 38724 95844 40348
rect 96012 38834 96068 41692
rect 96124 41186 96180 42812
rect 96348 41970 96404 43036
rect 97692 42756 97748 43596
rect 97692 42754 97860 42756
rect 97692 42702 97694 42754
rect 97746 42702 97860 42754
rect 97692 42700 97860 42702
rect 97692 42690 97748 42700
rect 97020 42644 97076 42654
rect 97020 42642 97300 42644
rect 97020 42590 97022 42642
rect 97074 42590 97300 42642
rect 97020 42588 97300 42590
rect 97020 42578 97076 42588
rect 97244 42194 97300 42588
rect 97244 42142 97246 42194
rect 97298 42142 97300 42194
rect 97244 42130 97300 42142
rect 96348 41918 96350 41970
rect 96402 41918 96404 41970
rect 96348 41906 96404 41918
rect 97468 41970 97524 41982
rect 97468 41918 97470 41970
rect 97522 41918 97524 41970
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 97132 41188 97188 41198
rect 96124 41134 96126 41186
rect 96178 41134 96180 41186
rect 96124 41122 96180 41134
rect 96908 41186 97188 41188
rect 96908 41134 97134 41186
rect 97186 41134 97188 41186
rect 96908 41132 97188 41134
rect 96796 41076 96852 41086
rect 96796 40982 96852 41020
rect 96348 40628 96404 40638
rect 96124 40516 96180 40526
rect 96124 40422 96180 40460
rect 96348 39058 96404 40572
rect 96908 40516 96964 41132
rect 97132 41122 97188 41132
rect 97356 41188 97412 41198
rect 97244 40516 97300 40526
rect 96908 40450 96964 40460
rect 97020 40514 97300 40516
rect 97020 40462 97246 40514
rect 97298 40462 97300 40514
rect 97020 40460 97300 40462
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 97020 39730 97076 40460
rect 97244 40450 97300 40460
rect 97020 39678 97022 39730
rect 97074 39678 97076 39730
rect 97020 39666 97076 39678
rect 96348 39006 96350 39058
rect 96402 39006 96404 39058
rect 96348 38994 96404 39006
rect 97132 39060 97188 39070
rect 97356 39060 97412 41132
rect 97468 40628 97524 41918
rect 97580 41188 97636 41198
rect 97580 41094 97636 41132
rect 97468 40562 97524 40572
rect 97132 39058 97412 39060
rect 97132 39006 97134 39058
rect 97186 39006 97412 39058
rect 97132 39004 97412 39006
rect 97468 40402 97524 40414
rect 97468 40350 97470 40402
rect 97522 40350 97524 40402
rect 97132 38994 97188 39004
rect 96012 38782 96014 38834
rect 96066 38782 96068 38834
rect 96012 38770 96068 38782
rect 96460 38836 96516 38846
rect 95788 38658 95844 38668
rect 95452 38546 95508 38556
rect 96236 38612 96292 38622
rect 95452 37940 95508 37950
rect 95452 37846 95508 37884
rect 95340 37326 95342 37378
rect 95394 37326 95396 37378
rect 93772 36642 93828 36652
rect 95228 36708 95284 36718
rect 95228 36614 95284 36652
rect 93212 36596 93268 36606
rect 93212 36502 93268 36540
rect 93772 36484 93828 36494
rect 93772 36390 93828 36428
rect 94332 36482 94388 36494
rect 94332 36430 94334 36482
rect 94386 36430 94388 36482
rect 92876 35186 92932 35196
rect 93660 34468 93716 34478
rect 93660 34354 93716 34412
rect 93660 34302 93662 34354
rect 93714 34302 93716 34354
rect 93660 34290 93716 34302
rect 93996 34468 94052 34478
rect 90188 33684 90244 33694
rect 90188 32562 90244 33628
rect 90188 32510 90190 32562
rect 90242 32510 90244 32562
rect 90188 32498 90244 32510
rect 90748 32674 90804 33964
rect 92204 34020 92260 34030
rect 92204 33926 92260 33964
rect 91644 33684 91700 33694
rect 91644 33458 91700 33628
rect 91644 33406 91646 33458
rect 91698 33406 91700 33458
rect 91644 33394 91700 33406
rect 92428 33348 92484 34076
rect 92764 34242 92820 34254
rect 92764 34190 92766 34242
rect 92818 34190 92820 34242
rect 92764 33684 92820 34190
rect 93100 34244 93156 34254
rect 93100 34150 93156 34188
rect 92764 33618 92820 33628
rect 92428 33254 92484 33292
rect 93996 33572 94052 34412
rect 94332 34356 94388 36430
rect 95340 36484 95396 37326
rect 95452 37266 95508 37278
rect 95452 37214 95454 37266
rect 95506 37214 95508 37266
rect 95452 36596 95508 37214
rect 95564 37268 95620 37278
rect 95564 36706 95620 37212
rect 96012 37268 96068 37278
rect 96012 37174 96068 37212
rect 95564 36654 95566 36706
rect 95618 36654 95620 36706
rect 95564 36642 95620 36654
rect 95452 36530 95508 36540
rect 95788 36596 95844 36606
rect 95340 36418 95396 36428
rect 95788 36370 95844 36540
rect 95788 36318 95790 36370
rect 95842 36318 95844 36370
rect 95788 36306 95844 36318
rect 96236 36596 96292 38556
rect 96348 37492 96404 37502
rect 96460 37492 96516 38780
rect 97468 38836 97524 40350
rect 97804 39620 97860 42700
rect 98028 41972 98084 41982
rect 98028 41878 98084 41916
rect 97916 41074 97972 41086
rect 97916 41022 97918 41074
rect 97970 41022 97972 41074
rect 97916 40628 97972 41022
rect 98028 40628 98084 40638
rect 97916 40626 98196 40628
rect 97916 40574 98030 40626
rect 98082 40574 98196 40626
rect 97916 40572 98196 40574
rect 98028 40562 98084 40572
rect 97580 39618 97972 39620
rect 97580 39566 97806 39618
rect 97858 39566 97972 39618
rect 97580 39564 97972 39566
rect 97580 39058 97636 39564
rect 97804 39554 97860 39564
rect 97580 39006 97582 39058
rect 97634 39006 97636 39058
rect 97580 38994 97636 39006
rect 97468 38770 97524 38780
rect 97020 38724 97076 38734
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 96348 37490 96516 37492
rect 96348 37438 96350 37490
rect 96402 37438 96516 37490
rect 96348 37436 96516 37438
rect 96348 37426 96404 37436
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 96908 36596 96964 36606
rect 96236 36594 96964 36596
rect 96236 36542 96910 36594
rect 96962 36542 96964 36594
rect 96236 36540 96964 36542
rect 96236 36370 96292 36540
rect 96908 36530 96964 36540
rect 96236 36318 96238 36370
rect 96290 36318 96292 36370
rect 94556 36260 94612 36270
rect 94556 36258 95172 36260
rect 94556 36206 94558 36258
rect 94610 36206 95172 36258
rect 94556 36204 95172 36206
rect 94556 36194 94612 36204
rect 94332 34290 94388 34300
rect 94444 35586 94500 35598
rect 94444 35534 94446 35586
rect 94498 35534 94500 35586
rect 94444 34914 94500 35534
rect 95116 35028 95172 36204
rect 96124 35252 96180 35262
rect 95116 34972 95396 35028
rect 94444 34862 94446 34914
rect 94498 34862 94500 34914
rect 93996 32788 94052 33516
rect 94332 34130 94388 34142
rect 94332 34078 94334 34130
rect 94386 34078 94388 34130
rect 94332 33124 94388 34078
rect 94444 33348 94500 34862
rect 95116 34804 95172 34814
rect 94556 34802 95172 34804
rect 94556 34750 95118 34802
rect 95170 34750 95172 34802
rect 94556 34748 95172 34750
rect 94556 34354 94612 34748
rect 95116 34738 95172 34748
rect 94556 34302 94558 34354
rect 94610 34302 94612 34354
rect 94556 34290 94612 34302
rect 95228 34356 95284 34366
rect 95228 34262 95284 34300
rect 95340 33458 95396 34972
rect 96124 34356 96180 35196
rect 95788 34242 95844 34254
rect 95788 34190 95790 34242
rect 95842 34190 95844 34242
rect 95340 33406 95342 33458
rect 95394 33406 95396 33458
rect 95340 33394 95396 33406
rect 95564 34132 95620 34142
rect 94556 33348 94612 33358
rect 94500 33346 94612 33348
rect 94500 33294 94558 33346
rect 94610 33294 94612 33346
rect 94500 33292 94612 33294
rect 94444 33216 94500 33292
rect 94556 33282 94612 33292
rect 94332 33068 95284 33124
rect 94108 32788 94164 32798
rect 93996 32786 94164 32788
rect 93996 32734 94110 32786
rect 94162 32734 94164 32786
rect 93996 32732 94164 32734
rect 94108 32722 94164 32732
rect 94668 32788 94724 32798
rect 94668 32694 94724 32732
rect 95228 32786 95284 33068
rect 95228 32734 95230 32786
rect 95282 32734 95284 32786
rect 95228 32722 95284 32734
rect 90748 32622 90750 32674
rect 90802 32622 90804 32674
rect 90748 31892 90804 32622
rect 90972 32564 91028 32574
rect 90972 32470 91028 32508
rect 91532 32564 91588 32574
rect 91532 32470 91588 32508
rect 95564 32562 95620 34076
rect 95788 33572 95844 34190
rect 96124 34242 96180 34300
rect 96124 34190 96126 34242
rect 96178 34190 96180 34242
rect 96124 34178 96180 34190
rect 95788 32674 95844 33516
rect 95788 32622 95790 32674
rect 95842 32622 95844 32674
rect 95788 32610 95844 32622
rect 96236 32788 96292 36318
rect 97020 35812 97076 38668
rect 97580 38162 97636 38174
rect 97580 38110 97582 38162
rect 97634 38110 97636 38162
rect 97580 37268 97636 38110
rect 97916 38164 97972 39564
rect 98028 38724 98084 38734
rect 98028 38630 98084 38668
rect 98140 38612 98196 40572
rect 98252 39732 98308 43652
rect 98252 39666 98308 39676
rect 98140 38546 98196 38556
rect 98028 38164 98084 38174
rect 97916 38162 98084 38164
rect 97916 38110 98030 38162
rect 98082 38110 98084 38162
rect 97916 38108 98084 38110
rect 98028 38098 98084 38108
rect 97580 37202 97636 37212
rect 97132 37154 97188 37166
rect 97132 37102 97134 37154
rect 97186 37102 97188 37154
rect 97132 36596 97188 37102
rect 97132 36530 97188 36540
rect 97132 35812 97188 35822
rect 96460 35810 97188 35812
rect 96460 35758 97134 35810
rect 97186 35758 97188 35810
rect 96460 35756 97188 35758
rect 96460 35698 96516 35756
rect 97132 35746 97188 35756
rect 96460 35646 96462 35698
rect 96514 35646 96516 35698
rect 96460 35634 96516 35646
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 97244 35026 97300 35038
rect 97244 34974 97246 35026
rect 97298 34974 97300 35026
rect 97132 34356 97188 34366
rect 97132 34262 97188 34300
rect 97244 34132 97300 34974
rect 97244 34066 97300 34076
rect 97468 34356 97524 34366
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 97468 33458 97524 34300
rect 97468 33406 97470 33458
rect 97522 33406 97524 33458
rect 97468 33394 97524 33406
rect 96236 32674 96292 32732
rect 96236 32622 96238 32674
rect 96290 32622 96292 32674
rect 96236 32610 96292 32622
rect 95564 32510 95566 32562
rect 95618 32510 95620 32562
rect 95564 32498 95620 32510
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 90748 31826 90804 31836
rect 90076 31614 90078 31666
rect 90130 31614 90132 31666
rect 90076 31602 90132 31614
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 95228 25394 95284 25406
rect 95228 25342 95230 25394
rect 95282 25342 95284 25394
rect 94892 25284 94948 25294
rect 94892 25190 94948 25228
rect 95228 25284 95284 25342
rect 95228 25218 95284 25228
rect 95788 25284 95844 25294
rect 95788 25190 95844 25228
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 93212 3444 93268 3454
rect 93436 3444 93492 3454
rect 93212 3442 93436 3444
rect 93212 3390 93214 3442
rect 93266 3390 93436 3442
rect 93212 3388 93436 3390
rect 93212 3378 93268 3388
rect 89628 3266 89684 3276
rect 82460 2930 82516 2940
rect 93436 800 93492 3388
rect 93996 3444 94052 3454
rect 93996 3350 94052 3388
rect 93660 3330 93716 3342
rect 93660 3278 93662 3330
rect 93714 3278 93716 3330
rect 93660 2884 93716 3278
rect 93660 2818 93716 2828
rect 6384 0 6496 800
rect 18816 0 18928 800
rect 31248 0 31360 800
rect 43680 0 43792 800
rect 56112 0 56224 800
rect 68544 0 68656 800
rect 80976 0 81088 800
rect 93408 0 93520 800
<< via2 >>
rect 4476 96458 4532 96460
rect 4476 96406 4478 96458
rect 4478 96406 4530 96458
rect 4530 96406 4532 96458
rect 4476 96404 4532 96406
rect 4580 96458 4636 96460
rect 4580 96406 4582 96458
rect 4582 96406 4634 96458
rect 4634 96406 4636 96458
rect 4580 96404 4636 96406
rect 4684 96458 4740 96460
rect 4684 96406 4686 96458
rect 4686 96406 4738 96458
rect 4738 96406 4740 96458
rect 4684 96404 4740 96406
rect 35196 96458 35252 96460
rect 35196 96406 35198 96458
rect 35198 96406 35250 96458
rect 35250 96406 35252 96458
rect 35196 96404 35252 96406
rect 35300 96458 35356 96460
rect 35300 96406 35302 96458
rect 35302 96406 35354 96458
rect 35354 96406 35356 96458
rect 35300 96404 35356 96406
rect 35404 96458 35460 96460
rect 35404 96406 35406 96458
rect 35406 96406 35458 96458
rect 35458 96406 35460 96458
rect 35404 96404 35460 96406
rect 65916 96458 65972 96460
rect 65916 96406 65918 96458
rect 65918 96406 65970 96458
rect 65970 96406 65972 96458
rect 65916 96404 65972 96406
rect 66020 96458 66076 96460
rect 66020 96406 66022 96458
rect 66022 96406 66074 96458
rect 66074 96406 66076 96458
rect 66020 96404 66076 96406
rect 66124 96458 66180 96460
rect 66124 96406 66126 96458
rect 66126 96406 66178 96458
rect 66178 96406 66180 96458
rect 66124 96404 66180 96406
rect 96636 96458 96692 96460
rect 96636 96406 96638 96458
rect 96638 96406 96690 96458
rect 96690 96406 96692 96458
rect 96636 96404 96692 96406
rect 96740 96458 96796 96460
rect 96740 96406 96742 96458
rect 96742 96406 96794 96458
rect 96794 96406 96796 96458
rect 96740 96404 96796 96406
rect 96844 96458 96900 96460
rect 96844 96406 96846 96458
rect 96846 96406 96898 96458
rect 96898 96406 96900 96458
rect 96844 96404 96900 96406
rect 93436 96124 93492 96180
rect 94332 96178 94388 96180
rect 94332 96126 94334 96178
rect 94334 96126 94386 96178
rect 94386 96126 94388 96178
rect 94332 96124 94388 96126
rect 7868 96066 7924 96068
rect 7868 96014 7870 96066
rect 7870 96014 7922 96066
rect 7922 96014 7924 96066
rect 7868 96012 7924 96014
rect 8316 96066 8372 96068
rect 8316 96014 8318 96066
rect 8318 96014 8370 96066
rect 8370 96014 8372 96066
rect 8316 96012 8372 96014
rect 20300 95788 20356 95844
rect 21308 95842 21364 95844
rect 21308 95790 21310 95842
rect 21310 95790 21362 95842
rect 21362 95790 21364 95842
rect 21308 95788 21364 95790
rect 27692 95788 27748 95844
rect 19836 95674 19892 95676
rect 19836 95622 19838 95674
rect 19838 95622 19890 95674
rect 19890 95622 19892 95674
rect 19836 95620 19892 95622
rect 19940 95674 19996 95676
rect 19940 95622 19942 95674
rect 19942 95622 19994 95674
rect 19994 95622 19996 95674
rect 19940 95620 19996 95622
rect 20044 95674 20100 95676
rect 20044 95622 20046 95674
rect 20046 95622 20098 95674
rect 20098 95622 20100 95674
rect 20044 95620 20100 95622
rect 4476 94890 4532 94892
rect 4476 94838 4478 94890
rect 4478 94838 4530 94890
rect 4530 94838 4532 94890
rect 4476 94836 4532 94838
rect 4580 94890 4636 94892
rect 4580 94838 4582 94890
rect 4582 94838 4634 94890
rect 4634 94838 4636 94890
rect 4580 94836 4636 94838
rect 4684 94890 4740 94892
rect 4684 94838 4686 94890
rect 4686 94838 4738 94890
rect 4738 94838 4740 94890
rect 4684 94836 4740 94838
rect 19836 94106 19892 94108
rect 19836 94054 19838 94106
rect 19838 94054 19890 94106
rect 19890 94054 19892 94106
rect 19836 94052 19892 94054
rect 19940 94106 19996 94108
rect 19940 94054 19942 94106
rect 19942 94054 19994 94106
rect 19994 94054 19996 94106
rect 19940 94052 19996 94054
rect 20044 94106 20100 94108
rect 20044 94054 20046 94106
rect 20046 94054 20098 94106
rect 20098 94054 20100 94106
rect 20044 94052 20100 94054
rect 4476 93322 4532 93324
rect 4476 93270 4478 93322
rect 4478 93270 4530 93322
rect 4530 93270 4532 93322
rect 4476 93268 4532 93270
rect 4580 93322 4636 93324
rect 4580 93270 4582 93322
rect 4582 93270 4634 93322
rect 4634 93270 4636 93322
rect 4580 93268 4636 93270
rect 4684 93322 4740 93324
rect 4684 93270 4686 93322
rect 4686 93270 4738 93322
rect 4738 93270 4740 93322
rect 4684 93268 4740 93270
rect 19836 92538 19892 92540
rect 19836 92486 19838 92538
rect 19838 92486 19890 92538
rect 19890 92486 19892 92538
rect 19836 92484 19892 92486
rect 19940 92538 19996 92540
rect 19940 92486 19942 92538
rect 19942 92486 19994 92538
rect 19994 92486 19996 92538
rect 19940 92484 19996 92486
rect 20044 92538 20100 92540
rect 20044 92486 20046 92538
rect 20046 92486 20098 92538
rect 20098 92486 20100 92538
rect 20044 92484 20100 92486
rect 4476 91754 4532 91756
rect 4476 91702 4478 91754
rect 4478 91702 4530 91754
rect 4530 91702 4532 91754
rect 4476 91700 4532 91702
rect 4580 91754 4636 91756
rect 4580 91702 4582 91754
rect 4582 91702 4634 91754
rect 4634 91702 4636 91754
rect 4580 91700 4636 91702
rect 4684 91754 4740 91756
rect 4684 91702 4686 91754
rect 4686 91702 4738 91754
rect 4738 91702 4740 91754
rect 4684 91700 4740 91702
rect 19836 90970 19892 90972
rect 19836 90918 19838 90970
rect 19838 90918 19890 90970
rect 19890 90918 19892 90970
rect 19836 90916 19892 90918
rect 19940 90970 19996 90972
rect 19940 90918 19942 90970
rect 19942 90918 19994 90970
rect 19994 90918 19996 90970
rect 19940 90916 19996 90918
rect 20044 90970 20100 90972
rect 20044 90918 20046 90970
rect 20046 90918 20098 90970
rect 20098 90918 20100 90970
rect 20044 90916 20100 90918
rect 4476 90186 4532 90188
rect 4476 90134 4478 90186
rect 4478 90134 4530 90186
rect 4530 90134 4532 90186
rect 4476 90132 4532 90134
rect 4580 90186 4636 90188
rect 4580 90134 4582 90186
rect 4582 90134 4634 90186
rect 4634 90134 4636 90186
rect 4580 90132 4636 90134
rect 4684 90186 4740 90188
rect 4684 90134 4686 90186
rect 4686 90134 4738 90186
rect 4738 90134 4740 90186
rect 4684 90132 4740 90134
rect 19836 89402 19892 89404
rect 19836 89350 19838 89402
rect 19838 89350 19890 89402
rect 19890 89350 19892 89402
rect 19836 89348 19892 89350
rect 19940 89402 19996 89404
rect 19940 89350 19942 89402
rect 19942 89350 19994 89402
rect 19994 89350 19996 89402
rect 19940 89348 19996 89350
rect 20044 89402 20100 89404
rect 20044 89350 20046 89402
rect 20046 89350 20098 89402
rect 20098 89350 20100 89402
rect 20044 89348 20100 89350
rect 4476 88618 4532 88620
rect 4476 88566 4478 88618
rect 4478 88566 4530 88618
rect 4530 88566 4532 88618
rect 4476 88564 4532 88566
rect 4580 88618 4636 88620
rect 4580 88566 4582 88618
rect 4582 88566 4634 88618
rect 4634 88566 4636 88618
rect 4580 88564 4636 88566
rect 4684 88618 4740 88620
rect 4684 88566 4686 88618
rect 4686 88566 4738 88618
rect 4738 88566 4740 88618
rect 4684 88564 4740 88566
rect 3276 88338 3332 88340
rect 3276 88286 3278 88338
rect 3278 88286 3330 88338
rect 3330 88286 3332 88338
rect 3276 88284 3332 88286
rect 12572 88284 12628 88340
rect 1708 87442 1764 87444
rect 1708 87390 1710 87442
rect 1710 87390 1762 87442
rect 1762 87390 1764 87442
rect 1708 87388 1764 87390
rect 4476 87050 4532 87052
rect 4476 86998 4478 87050
rect 4478 86998 4530 87050
rect 4530 86998 4532 87050
rect 4476 86996 4532 86998
rect 4580 87050 4636 87052
rect 4580 86998 4582 87050
rect 4582 86998 4634 87050
rect 4634 86998 4636 87050
rect 4580 86996 4636 86998
rect 4684 87050 4740 87052
rect 4684 86998 4686 87050
rect 4686 86998 4738 87050
rect 4738 86998 4740 87050
rect 4684 86996 4740 86998
rect 4476 85482 4532 85484
rect 4476 85430 4478 85482
rect 4478 85430 4530 85482
rect 4530 85430 4532 85482
rect 4476 85428 4532 85430
rect 4580 85482 4636 85484
rect 4580 85430 4582 85482
rect 4582 85430 4634 85482
rect 4634 85430 4636 85482
rect 4580 85428 4636 85430
rect 4684 85482 4740 85484
rect 4684 85430 4686 85482
rect 4686 85430 4738 85482
rect 4738 85430 4740 85482
rect 4684 85428 4740 85430
rect 4476 83914 4532 83916
rect 4476 83862 4478 83914
rect 4478 83862 4530 83914
rect 4530 83862 4532 83914
rect 4476 83860 4532 83862
rect 4580 83914 4636 83916
rect 4580 83862 4582 83914
rect 4582 83862 4634 83914
rect 4634 83862 4636 83914
rect 4580 83860 4636 83862
rect 4684 83914 4740 83916
rect 4684 83862 4686 83914
rect 4686 83862 4738 83914
rect 4738 83862 4740 83914
rect 4684 83860 4740 83862
rect 4476 82346 4532 82348
rect 4476 82294 4478 82346
rect 4478 82294 4530 82346
rect 4530 82294 4532 82346
rect 4476 82292 4532 82294
rect 4580 82346 4636 82348
rect 4580 82294 4582 82346
rect 4582 82294 4634 82346
rect 4634 82294 4636 82346
rect 4580 82292 4636 82294
rect 4684 82346 4740 82348
rect 4684 82294 4686 82346
rect 4686 82294 4738 82346
rect 4738 82294 4740 82346
rect 4684 82292 4740 82294
rect 4476 80778 4532 80780
rect 4476 80726 4478 80778
rect 4478 80726 4530 80778
rect 4530 80726 4532 80778
rect 4476 80724 4532 80726
rect 4580 80778 4636 80780
rect 4580 80726 4582 80778
rect 4582 80726 4634 80778
rect 4634 80726 4636 80778
rect 4580 80724 4636 80726
rect 4684 80778 4740 80780
rect 4684 80726 4686 80778
rect 4686 80726 4738 80778
rect 4738 80726 4740 80778
rect 4684 80724 4740 80726
rect 4476 79210 4532 79212
rect 4476 79158 4478 79210
rect 4478 79158 4530 79210
rect 4530 79158 4532 79210
rect 4476 79156 4532 79158
rect 4580 79210 4636 79212
rect 4580 79158 4582 79210
rect 4582 79158 4634 79210
rect 4634 79158 4636 79210
rect 4580 79156 4636 79158
rect 4684 79210 4740 79212
rect 4684 79158 4686 79210
rect 4686 79158 4738 79210
rect 4738 79158 4740 79210
rect 4684 79156 4740 79158
rect 4476 77642 4532 77644
rect 4476 77590 4478 77642
rect 4478 77590 4530 77642
rect 4530 77590 4532 77642
rect 4476 77588 4532 77590
rect 4580 77642 4636 77644
rect 4580 77590 4582 77642
rect 4582 77590 4634 77642
rect 4634 77590 4636 77642
rect 4580 77588 4636 77590
rect 4684 77642 4740 77644
rect 4684 77590 4686 77642
rect 4686 77590 4738 77642
rect 4738 77590 4740 77642
rect 4684 77588 4740 77590
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 19836 87834 19892 87836
rect 19836 87782 19838 87834
rect 19838 87782 19890 87834
rect 19890 87782 19892 87834
rect 19836 87780 19892 87782
rect 19940 87834 19996 87836
rect 19940 87782 19942 87834
rect 19942 87782 19994 87834
rect 19994 87782 19996 87834
rect 19940 87780 19996 87782
rect 20044 87834 20100 87836
rect 20044 87782 20046 87834
rect 20046 87782 20098 87834
rect 20098 87782 20100 87834
rect 20044 87780 20100 87782
rect 19836 86266 19892 86268
rect 19836 86214 19838 86266
rect 19838 86214 19890 86266
rect 19890 86214 19892 86266
rect 19836 86212 19892 86214
rect 19940 86266 19996 86268
rect 19940 86214 19942 86266
rect 19942 86214 19994 86266
rect 19994 86214 19996 86266
rect 19940 86212 19996 86214
rect 20044 86266 20100 86268
rect 20044 86214 20046 86266
rect 20046 86214 20098 86266
rect 20098 86214 20100 86266
rect 20044 86212 20100 86214
rect 19836 84698 19892 84700
rect 19836 84646 19838 84698
rect 19838 84646 19890 84698
rect 19890 84646 19892 84698
rect 19836 84644 19892 84646
rect 19940 84698 19996 84700
rect 19940 84646 19942 84698
rect 19942 84646 19994 84698
rect 19994 84646 19996 84698
rect 19940 84644 19996 84646
rect 20044 84698 20100 84700
rect 20044 84646 20046 84698
rect 20046 84646 20098 84698
rect 20098 84646 20100 84698
rect 20044 84644 20100 84646
rect 19836 83130 19892 83132
rect 19836 83078 19838 83130
rect 19838 83078 19890 83130
rect 19890 83078 19892 83130
rect 19836 83076 19892 83078
rect 19940 83130 19996 83132
rect 19940 83078 19942 83130
rect 19942 83078 19994 83130
rect 19994 83078 19996 83130
rect 19940 83076 19996 83078
rect 20044 83130 20100 83132
rect 20044 83078 20046 83130
rect 20046 83078 20098 83130
rect 20098 83078 20100 83130
rect 20044 83076 20100 83078
rect 19836 81562 19892 81564
rect 19836 81510 19838 81562
rect 19838 81510 19890 81562
rect 19890 81510 19892 81562
rect 19836 81508 19892 81510
rect 19940 81562 19996 81564
rect 19940 81510 19942 81562
rect 19942 81510 19994 81562
rect 19994 81510 19996 81562
rect 19940 81508 19996 81510
rect 20044 81562 20100 81564
rect 20044 81510 20046 81562
rect 20046 81510 20098 81562
rect 20098 81510 20100 81562
rect 20044 81508 20100 81510
rect 19836 79994 19892 79996
rect 19836 79942 19838 79994
rect 19838 79942 19890 79994
rect 19890 79942 19892 79994
rect 19836 79940 19892 79942
rect 19940 79994 19996 79996
rect 19940 79942 19942 79994
rect 19942 79942 19994 79994
rect 19994 79942 19996 79994
rect 19940 79940 19996 79942
rect 20044 79994 20100 79996
rect 20044 79942 20046 79994
rect 20046 79942 20098 79994
rect 20098 79942 20100 79994
rect 20044 79940 20100 79942
rect 19836 78426 19892 78428
rect 19836 78374 19838 78426
rect 19838 78374 19890 78426
rect 19890 78374 19892 78426
rect 19836 78372 19892 78374
rect 19940 78426 19996 78428
rect 19940 78374 19942 78426
rect 19942 78374 19994 78426
rect 19994 78374 19996 78426
rect 19940 78372 19996 78374
rect 20044 78426 20100 78428
rect 20044 78374 20046 78426
rect 20046 78374 20098 78426
rect 20098 78374 20100 78426
rect 20044 78372 20100 78374
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 27692 64764 27748 64820
rect 47964 96012 48020 96068
rect 35196 94890 35252 94892
rect 35196 94838 35198 94890
rect 35198 94838 35250 94890
rect 35250 94838 35252 94890
rect 35196 94836 35252 94838
rect 35300 94890 35356 94892
rect 35300 94838 35302 94890
rect 35302 94838 35354 94890
rect 35354 94838 35356 94890
rect 35300 94836 35356 94838
rect 35404 94890 35460 94892
rect 35404 94838 35406 94890
rect 35406 94838 35458 94890
rect 35458 94838 35460 94890
rect 35404 94836 35460 94838
rect 35196 93322 35252 93324
rect 35196 93270 35198 93322
rect 35198 93270 35250 93322
rect 35250 93270 35252 93322
rect 35196 93268 35252 93270
rect 35300 93322 35356 93324
rect 35300 93270 35302 93322
rect 35302 93270 35354 93322
rect 35354 93270 35356 93322
rect 35300 93268 35356 93270
rect 35404 93322 35460 93324
rect 35404 93270 35406 93322
rect 35406 93270 35458 93322
rect 35458 93270 35460 93322
rect 35404 93268 35460 93270
rect 35196 91754 35252 91756
rect 35196 91702 35198 91754
rect 35198 91702 35250 91754
rect 35250 91702 35252 91754
rect 35196 91700 35252 91702
rect 35300 91754 35356 91756
rect 35300 91702 35302 91754
rect 35302 91702 35354 91754
rect 35354 91702 35356 91754
rect 35300 91700 35356 91702
rect 35404 91754 35460 91756
rect 35404 91702 35406 91754
rect 35406 91702 35458 91754
rect 35458 91702 35460 91754
rect 35404 91700 35460 91702
rect 35196 90186 35252 90188
rect 35196 90134 35198 90186
rect 35198 90134 35250 90186
rect 35250 90134 35252 90186
rect 35196 90132 35252 90134
rect 35300 90186 35356 90188
rect 35300 90134 35302 90186
rect 35302 90134 35354 90186
rect 35354 90134 35356 90186
rect 35300 90132 35356 90134
rect 35404 90186 35460 90188
rect 35404 90134 35406 90186
rect 35406 90134 35458 90186
rect 35458 90134 35460 90186
rect 35404 90132 35460 90134
rect 35196 88618 35252 88620
rect 35196 88566 35198 88618
rect 35198 88566 35250 88618
rect 35250 88566 35252 88618
rect 35196 88564 35252 88566
rect 35300 88618 35356 88620
rect 35300 88566 35302 88618
rect 35302 88566 35354 88618
rect 35354 88566 35356 88618
rect 35300 88564 35356 88566
rect 35404 88618 35460 88620
rect 35404 88566 35406 88618
rect 35406 88566 35458 88618
rect 35458 88566 35460 88618
rect 35404 88564 35460 88566
rect 35196 87050 35252 87052
rect 35196 86998 35198 87050
rect 35198 86998 35250 87050
rect 35250 86998 35252 87050
rect 35196 86996 35252 86998
rect 35300 87050 35356 87052
rect 35300 86998 35302 87050
rect 35302 86998 35354 87050
rect 35354 86998 35356 87050
rect 35300 86996 35356 86998
rect 35404 87050 35460 87052
rect 35404 86998 35406 87050
rect 35406 86998 35458 87050
rect 35458 86998 35460 87050
rect 35404 86996 35460 86998
rect 35196 85482 35252 85484
rect 35196 85430 35198 85482
rect 35198 85430 35250 85482
rect 35250 85430 35252 85482
rect 35196 85428 35252 85430
rect 35300 85482 35356 85484
rect 35300 85430 35302 85482
rect 35302 85430 35354 85482
rect 35354 85430 35356 85482
rect 35300 85428 35356 85430
rect 35404 85482 35460 85484
rect 35404 85430 35406 85482
rect 35406 85430 35458 85482
rect 35458 85430 35460 85482
rect 35404 85428 35460 85430
rect 35196 83914 35252 83916
rect 35196 83862 35198 83914
rect 35198 83862 35250 83914
rect 35250 83862 35252 83914
rect 35196 83860 35252 83862
rect 35300 83914 35356 83916
rect 35300 83862 35302 83914
rect 35302 83862 35354 83914
rect 35354 83862 35356 83914
rect 35300 83860 35356 83862
rect 35404 83914 35460 83916
rect 35404 83862 35406 83914
rect 35406 83862 35458 83914
rect 35458 83862 35460 83914
rect 35404 83860 35460 83862
rect 35196 82346 35252 82348
rect 35196 82294 35198 82346
rect 35198 82294 35250 82346
rect 35250 82294 35252 82346
rect 35196 82292 35252 82294
rect 35300 82346 35356 82348
rect 35300 82294 35302 82346
rect 35302 82294 35354 82346
rect 35354 82294 35356 82346
rect 35300 82292 35356 82294
rect 35404 82346 35460 82348
rect 35404 82294 35406 82346
rect 35406 82294 35458 82346
rect 35458 82294 35460 82346
rect 35404 82292 35460 82294
rect 35196 80778 35252 80780
rect 35196 80726 35198 80778
rect 35198 80726 35250 80778
rect 35250 80726 35252 80778
rect 35196 80724 35252 80726
rect 35300 80778 35356 80780
rect 35300 80726 35302 80778
rect 35302 80726 35354 80778
rect 35354 80726 35356 80778
rect 35300 80724 35356 80726
rect 35404 80778 35460 80780
rect 35404 80726 35406 80778
rect 35406 80726 35458 80778
rect 35458 80726 35460 80778
rect 35404 80724 35460 80726
rect 35196 79210 35252 79212
rect 35196 79158 35198 79210
rect 35198 79158 35250 79210
rect 35250 79158 35252 79210
rect 35196 79156 35252 79158
rect 35300 79210 35356 79212
rect 35300 79158 35302 79210
rect 35302 79158 35354 79210
rect 35354 79158 35356 79210
rect 35300 79156 35356 79158
rect 35404 79210 35460 79212
rect 35404 79158 35406 79210
rect 35406 79158 35458 79210
rect 35458 79158 35460 79210
rect 35404 79156 35460 79158
rect 35196 77642 35252 77644
rect 35196 77590 35198 77642
rect 35198 77590 35250 77642
rect 35250 77590 35252 77642
rect 35196 77588 35252 77590
rect 35300 77642 35356 77644
rect 35300 77590 35302 77642
rect 35302 77590 35354 77642
rect 35354 77590 35356 77642
rect 35300 77588 35356 77590
rect 35404 77642 35460 77644
rect 35404 77590 35406 77642
rect 35406 77590 35458 77642
rect 35458 77590 35460 77642
rect 35404 77588 35460 77590
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 47852 68908 47908 68964
rect 45948 68684 46004 68740
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 32172 64652 32228 64708
rect 46956 64652 47012 64708
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 12572 63644 12628 63700
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 46956 63532 47012 63588
rect 35404 63476 35460 63478
rect 50556 95674 50612 95676
rect 50556 95622 50558 95674
rect 50558 95622 50610 95674
rect 50610 95622 50612 95674
rect 50556 95620 50612 95622
rect 50660 95674 50716 95676
rect 50660 95622 50662 95674
rect 50662 95622 50714 95674
rect 50714 95622 50716 95674
rect 50660 95620 50716 95622
rect 50764 95674 50820 95676
rect 50764 95622 50766 95674
rect 50766 95622 50818 95674
rect 50818 95622 50820 95674
rect 50764 95620 50820 95622
rect 50556 94106 50612 94108
rect 50556 94054 50558 94106
rect 50558 94054 50610 94106
rect 50610 94054 50612 94106
rect 50556 94052 50612 94054
rect 50660 94106 50716 94108
rect 50660 94054 50662 94106
rect 50662 94054 50714 94106
rect 50714 94054 50716 94106
rect 50660 94052 50716 94054
rect 50764 94106 50820 94108
rect 50764 94054 50766 94106
rect 50766 94054 50818 94106
rect 50818 94054 50820 94106
rect 50764 94052 50820 94054
rect 50556 92538 50612 92540
rect 50556 92486 50558 92538
rect 50558 92486 50610 92538
rect 50610 92486 50612 92538
rect 50556 92484 50612 92486
rect 50660 92538 50716 92540
rect 50660 92486 50662 92538
rect 50662 92486 50714 92538
rect 50714 92486 50716 92538
rect 50660 92484 50716 92486
rect 50764 92538 50820 92540
rect 50764 92486 50766 92538
rect 50766 92486 50818 92538
rect 50818 92486 50820 92538
rect 50764 92484 50820 92486
rect 50556 90970 50612 90972
rect 50556 90918 50558 90970
rect 50558 90918 50610 90970
rect 50610 90918 50612 90970
rect 50556 90916 50612 90918
rect 50660 90970 50716 90972
rect 50660 90918 50662 90970
rect 50662 90918 50714 90970
rect 50714 90918 50716 90970
rect 50660 90916 50716 90918
rect 50764 90970 50820 90972
rect 50764 90918 50766 90970
rect 50766 90918 50818 90970
rect 50818 90918 50820 90970
rect 50764 90916 50820 90918
rect 50556 89402 50612 89404
rect 50556 89350 50558 89402
rect 50558 89350 50610 89402
rect 50610 89350 50612 89402
rect 50556 89348 50612 89350
rect 50660 89402 50716 89404
rect 50660 89350 50662 89402
rect 50662 89350 50714 89402
rect 50714 89350 50716 89402
rect 50660 89348 50716 89350
rect 50764 89402 50820 89404
rect 50764 89350 50766 89402
rect 50766 89350 50818 89402
rect 50818 89350 50820 89402
rect 50764 89348 50820 89350
rect 50556 87834 50612 87836
rect 50556 87782 50558 87834
rect 50558 87782 50610 87834
rect 50610 87782 50612 87834
rect 50556 87780 50612 87782
rect 50660 87834 50716 87836
rect 50660 87782 50662 87834
rect 50662 87782 50714 87834
rect 50714 87782 50716 87834
rect 50660 87780 50716 87782
rect 50764 87834 50820 87836
rect 50764 87782 50766 87834
rect 50766 87782 50818 87834
rect 50818 87782 50820 87834
rect 50764 87780 50820 87782
rect 54236 87276 54292 87332
rect 53564 87218 53620 87220
rect 53564 87166 53566 87218
rect 53566 87166 53618 87218
rect 53618 87166 53620 87218
rect 53564 87164 53620 87166
rect 50556 86266 50612 86268
rect 50556 86214 50558 86266
rect 50558 86214 50610 86266
rect 50610 86214 50612 86266
rect 50556 86212 50612 86214
rect 50660 86266 50716 86268
rect 50660 86214 50662 86266
rect 50662 86214 50714 86266
rect 50714 86214 50716 86266
rect 50660 86212 50716 86214
rect 50764 86266 50820 86268
rect 50764 86214 50766 86266
rect 50766 86214 50818 86266
rect 50818 86214 50820 86266
rect 50764 86212 50820 86214
rect 50556 84698 50612 84700
rect 50556 84646 50558 84698
rect 50558 84646 50610 84698
rect 50610 84646 50612 84698
rect 50556 84644 50612 84646
rect 50660 84698 50716 84700
rect 50660 84646 50662 84698
rect 50662 84646 50714 84698
rect 50714 84646 50716 84698
rect 50660 84644 50716 84646
rect 50764 84698 50820 84700
rect 50764 84646 50766 84698
rect 50766 84646 50818 84698
rect 50818 84646 50820 84698
rect 50764 84644 50820 84646
rect 54012 85932 54068 85988
rect 54796 87276 54852 87332
rect 55020 87330 55076 87332
rect 55020 87278 55022 87330
rect 55022 87278 55074 87330
rect 55074 87278 55076 87330
rect 55020 87276 55076 87278
rect 53788 84866 53844 84868
rect 53788 84814 53790 84866
rect 53790 84814 53842 84866
rect 53842 84814 53844 84866
rect 53788 84812 53844 84814
rect 50556 83130 50612 83132
rect 50556 83078 50558 83130
rect 50558 83078 50610 83130
rect 50610 83078 50612 83130
rect 50556 83076 50612 83078
rect 50660 83130 50716 83132
rect 50660 83078 50662 83130
rect 50662 83078 50714 83130
rect 50714 83078 50716 83130
rect 50660 83076 50716 83078
rect 50764 83130 50820 83132
rect 50764 83078 50766 83130
rect 50766 83078 50818 83130
rect 50818 83078 50820 83130
rect 50764 83076 50820 83078
rect 50556 81562 50612 81564
rect 50556 81510 50558 81562
rect 50558 81510 50610 81562
rect 50610 81510 50612 81562
rect 50556 81508 50612 81510
rect 50660 81562 50716 81564
rect 50660 81510 50662 81562
rect 50662 81510 50714 81562
rect 50714 81510 50716 81562
rect 50660 81508 50716 81510
rect 50764 81562 50820 81564
rect 50764 81510 50766 81562
rect 50766 81510 50818 81562
rect 50818 81510 50820 81562
rect 50764 81508 50820 81510
rect 49756 81116 49812 81172
rect 49308 78706 49364 78708
rect 49308 78654 49310 78706
rect 49310 78654 49362 78706
rect 49362 78654 49364 78706
rect 49308 78652 49364 78654
rect 49756 78594 49812 78596
rect 49756 78542 49758 78594
rect 49758 78542 49810 78594
rect 49810 78542 49812 78594
rect 49756 78540 49812 78542
rect 48860 78258 48916 78260
rect 48860 78206 48862 78258
rect 48862 78206 48914 78258
rect 48914 78206 48916 78258
rect 48860 78204 48916 78206
rect 49644 78204 49700 78260
rect 48300 78146 48356 78148
rect 48300 78094 48302 78146
rect 48302 78094 48354 78146
rect 48354 78094 48356 78146
rect 48300 78092 48356 78094
rect 50316 81282 50372 81284
rect 50316 81230 50318 81282
rect 50318 81230 50370 81282
rect 50370 81230 50372 81282
rect 50316 81228 50372 81230
rect 50556 79994 50612 79996
rect 50556 79942 50558 79994
rect 50558 79942 50610 79994
rect 50610 79942 50612 79994
rect 50556 79940 50612 79942
rect 50660 79994 50716 79996
rect 50660 79942 50662 79994
rect 50662 79942 50714 79994
rect 50714 79942 50716 79994
rect 50660 79940 50716 79942
rect 50764 79994 50820 79996
rect 50764 79942 50766 79994
rect 50766 79942 50818 79994
rect 50818 79942 50820 79994
rect 50764 79940 50820 79942
rect 50204 78764 50260 78820
rect 50092 78652 50148 78708
rect 49756 78146 49812 78148
rect 49756 78094 49758 78146
rect 49758 78094 49810 78146
rect 49810 78094 49812 78146
rect 49756 78092 49812 78094
rect 50764 78706 50820 78708
rect 50764 78654 50766 78706
rect 50766 78654 50818 78706
rect 50818 78654 50820 78706
rect 50764 78652 50820 78654
rect 50204 78594 50260 78596
rect 50204 78542 50206 78594
rect 50206 78542 50258 78594
rect 50258 78542 50260 78594
rect 50204 78540 50260 78542
rect 50556 78426 50612 78428
rect 50556 78374 50558 78426
rect 50558 78374 50610 78426
rect 50610 78374 50612 78426
rect 50556 78372 50612 78374
rect 50660 78426 50716 78428
rect 50660 78374 50662 78426
rect 50662 78374 50714 78426
rect 50714 78374 50716 78426
rect 50660 78372 50716 78374
rect 50764 78426 50820 78428
rect 50764 78374 50766 78426
rect 50766 78374 50818 78426
rect 50818 78374 50820 78426
rect 50764 78372 50820 78374
rect 50428 78204 50484 78260
rect 50092 77308 50148 77364
rect 50316 78092 50372 78148
rect 49868 76972 49924 77028
rect 54684 86044 54740 86100
rect 54460 84812 54516 84868
rect 56028 87164 56084 87220
rect 56476 86716 56532 86772
rect 57484 87164 57540 87220
rect 70028 95788 70084 95844
rect 70476 95842 70532 95844
rect 70476 95790 70478 95842
rect 70478 95790 70530 95842
rect 70530 95790 70532 95842
rect 70476 95788 70532 95790
rect 77980 95788 78036 95844
rect 65916 94890 65972 94892
rect 65916 94838 65918 94890
rect 65918 94838 65970 94890
rect 65970 94838 65972 94890
rect 65916 94836 65972 94838
rect 66020 94890 66076 94892
rect 66020 94838 66022 94890
rect 66022 94838 66074 94890
rect 66074 94838 66076 94890
rect 66020 94836 66076 94838
rect 66124 94890 66180 94892
rect 66124 94838 66126 94890
rect 66126 94838 66178 94890
rect 66178 94838 66180 94890
rect 66124 94836 66180 94838
rect 65916 93322 65972 93324
rect 65916 93270 65918 93322
rect 65918 93270 65970 93322
rect 65970 93270 65972 93322
rect 65916 93268 65972 93270
rect 66020 93322 66076 93324
rect 66020 93270 66022 93322
rect 66022 93270 66074 93322
rect 66074 93270 66076 93322
rect 66020 93268 66076 93270
rect 66124 93322 66180 93324
rect 66124 93270 66126 93322
rect 66126 93270 66178 93322
rect 66178 93270 66180 93322
rect 66124 93268 66180 93270
rect 65916 91754 65972 91756
rect 65916 91702 65918 91754
rect 65918 91702 65970 91754
rect 65970 91702 65972 91754
rect 65916 91700 65972 91702
rect 66020 91754 66076 91756
rect 66020 91702 66022 91754
rect 66022 91702 66074 91754
rect 66074 91702 66076 91754
rect 66020 91700 66076 91702
rect 66124 91754 66180 91756
rect 66124 91702 66126 91754
rect 66126 91702 66178 91754
rect 66178 91702 66180 91754
rect 66124 91700 66180 91702
rect 93100 96066 93156 96068
rect 93100 96014 93102 96066
rect 93102 96014 93154 96066
rect 93154 96014 93156 96066
rect 93100 96012 93156 96014
rect 93884 96066 93940 96068
rect 93884 96014 93886 96066
rect 93886 96014 93938 96066
rect 93938 96014 93940 96066
rect 93884 96012 93940 96014
rect 97468 96012 97524 96068
rect 81276 95674 81332 95676
rect 81276 95622 81278 95674
rect 81278 95622 81330 95674
rect 81330 95622 81332 95674
rect 81276 95620 81332 95622
rect 81380 95674 81436 95676
rect 81380 95622 81382 95674
rect 81382 95622 81434 95674
rect 81434 95622 81436 95674
rect 81380 95620 81436 95622
rect 81484 95674 81540 95676
rect 81484 95622 81486 95674
rect 81486 95622 81538 95674
rect 81538 95622 81540 95674
rect 81484 95620 81540 95622
rect 81276 94106 81332 94108
rect 81276 94054 81278 94106
rect 81278 94054 81330 94106
rect 81330 94054 81332 94106
rect 81276 94052 81332 94054
rect 81380 94106 81436 94108
rect 81380 94054 81382 94106
rect 81382 94054 81434 94106
rect 81434 94054 81436 94106
rect 81380 94052 81436 94054
rect 81484 94106 81540 94108
rect 81484 94054 81486 94106
rect 81486 94054 81538 94106
rect 81538 94054 81540 94106
rect 81484 94052 81540 94054
rect 81276 92538 81332 92540
rect 81276 92486 81278 92538
rect 81278 92486 81330 92538
rect 81330 92486 81332 92538
rect 81276 92484 81332 92486
rect 81380 92538 81436 92540
rect 81380 92486 81382 92538
rect 81382 92486 81434 92538
rect 81434 92486 81436 92538
rect 81380 92484 81436 92486
rect 81484 92538 81540 92540
rect 81484 92486 81486 92538
rect 81486 92486 81538 92538
rect 81538 92486 81540 92538
rect 81484 92484 81540 92486
rect 81276 90970 81332 90972
rect 81276 90918 81278 90970
rect 81278 90918 81330 90970
rect 81330 90918 81332 90970
rect 81276 90916 81332 90918
rect 81380 90970 81436 90972
rect 81380 90918 81382 90970
rect 81382 90918 81434 90970
rect 81434 90918 81436 90970
rect 81380 90916 81436 90918
rect 81484 90970 81540 90972
rect 81484 90918 81486 90970
rect 81486 90918 81538 90970
rect 81538 90918 81540 90970
rect 81484 90916 81540 90918
rect 65916 90186 65972 90188
rect 65916 90134 65918 90186
rect 65918 90134 65970 90186
rect 65970 90134 65972 90186
rect 65916 90132 65972 90134
rect 66020 90186 66076 90188
rect 66020 90134 66022 90186
rect 66022 90134 66074 90186
rect 66074 90134 66076 90186
rect 66020 90132 66076 90134
rect 66124 90186 66180 90188
rect 66124 90134 66126 90186
rect 66126 90134 66178 90186
rect 66178 90134 66180 90186
rect 66124 90132 66180 90134
rect 59052 87836 59108 87892
rect 59612 87836 59668 87892
rect 60284 87836 60340 87892
rect 57596 86940 57652 86996
rect 57820 87164 57876 87220
rect 57596 86716 57652 86772
rect 55692 85932 55748 85988
rect 56476 86044 56532 86100
rect 55804 85762 55860 85764
rect 55804 85710 55806 85762
rect 55806 85710 55858 85762
rect 55858 85710 55860 85762
rect 55804 85708 55860 85710
rect 53228 83580 53284 83636
rect 52444 83244 52500 83300
rect 52220 82684 52276 82740
rect 51212 81116 51268 81172
rect 51660 81170 51716 81172
rect 51660 81118 51662 81170
rect 51662 81118 51714 81170
rect 51714 81118 51716 81170
rect 51660 81116 51716 81118
rect 51100 80892 51156 80948
rect 52108 78818 52164 78820
rect 52108 78766 52110 78818
rect 52110 78766 52162 78818
rect 52162 78766 52164 78818
rect 52108 78764 52164 78766
rect 50988 78594 51044 78596
rect 50988 78542 50990 78594
rect 50990 78542 51042 78594
rect 51042 78542 51044 78594
rect 50988 78540 51044 78542
rect 50540 77980 50596 78036
rect 51324 78146 51380 78148
rect 51324 78094 51326 78146
rect 51326 78094 51378 78146
rect 51378 78094 51380 78146
rect 51324 78092 51380 78094
rect 51212 77868 51268 77924
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50204 74226 50260 74228
rect 50204 74174 50206 74226
rect 50206 74174 50258 74226
rect 50258 74174 50260 74226
rect 50204 74172 50260 74174
rect 49756 71932 49812 71988
rect 48188 70866 48244 70868
rect 48188 70814 48190 70866
rect 48190 70814 48242 70866
rect 48242 70814 48244 70866
rect 48188 70812 48244 70814
rect 47964 63196 48020 63252
rect 48076 70700 48132 70756
rect 2156 62748 2212 62804
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 1820 62466 1876 62468
rect 1820 62414 1822 62466
rect 1822 62414 1874 62466
rect 1874 62414 1876 62466
rect 1820 62412 1876 62414
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 49532 70866 49588 70868
rect 49532 70814 49534 70866
rect 49534 70814 49586 70866
rect 49586 70814 49588 70866
rect 49532 70812 49588 70814
rect 48972 69356 49028 69412
rect 49532 69410 49588 69412
rect 49532 69358 49534 69410
rect 49534 69358 49586 69410
rect 49586 69358 49588 69410
rect 49532 69356 49588 69358
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50764 75010 50820 75012
rect 50764 74958 50766 75010
rect 50766 74958 50818 75010
rect 50818 74958 50820 75010
rect 50764 74956 50820 74958
rect 50652 74172 50708 74228
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 52668 82066 52724 82068
rect 52668 82014 52670 82066
rect 52670 82014 52722 82066
rect 52722 82014 52724 82066
rect 52668 82012 52724 82014
rect 52892 82738 52948 82740
rect 52892 82686 52894 82738
rect 52894 82686 52946 82738
rect 52946 82686 52948 82738
rect 52892 82684 52948 82686
rect 52780 81900 52836 81956
rect 52332 79772 52388 79828
rect 52892 79826 52948 79828
rect 52892 79774 52894 79826
rect 52894 79774 52946 79826
rect 52946 79774 52948 79826
rect 52892 79772 52948 79774
rect 53676 83580 53732 83636
rect 56588 85148 56644 85204
rect 56700 85932 56756 85988
rect 54460 83580 54516 83636
rect 53340 81900 53396 81956
rect 53340 81116 53396 81172
rect 54124 83298 54180 83300
rect 54124 83246 54126 83298
rect 54126 83246 54178 83298
rect 54178 83246 54180 83298
rect 54124 83244 54180 83246
rect 53564 82012 53620 82068
rect 54124 82236 54180 82292
rect 54124 81954 54180 81956
rect 54124 81902 54126 81954
rect 54126 81902 54178 81954
rect 54178 81902 54180 81954
rect 54124 81900 54180 81902
rect 53452 80892 53508 80948
rect 54012 81228 54068 81284
rect 53228 80108 53284 80164
rect 55804 84140 55860 84196
rect 56476 84140 56532 84196
rect 54908 82236 54964 82292
rect 55020 81676 55076 81732
rect 54236 80498 54292 80500
rect 54236 80446 54238 80498
rect 54238 80446 54290 80498
rect 54290 80446 54292 80498
rect 54236 80444 54292 80446
rect 53676 78988 53732 79044
rect 53340 78818 53396 78820
rect 53340 78766 53342 78818
rect 53342 78766 53394 78818
rect 53394 78766 53396 78818
rect 53340 78764 53396 78766
rect 52332 78594 52388 78596
rect 52332 78542 52334 78594
rect 52334 78542 52386 78594
rect 52386 78542 52388 78594
rect 52332 78540 52388 78542
rect 51660 77084 51716 77140
rect 51772 77980 51828 78036
rect 51660 75180 51716 75236
rect 51884 74956 51940 75012
rect 51996 77308 52052 77364
rect 54908 80444 54964 80500
rect 55020 80892 55076 80948
rect 54572 79714 54628 79716
rect 54572 79662 54574 79714
rect 54574 79662 54626 79714
rect 54626 79662 54628 79714
rect 54572 79660 54628 79662
rect 54684 79602 54740 79604
rect 54684 79550 54686 79602
rect 54686 79550 54738 79602
rect 54738 79550 54740 79602
rect 54684 79548 54740 79550
rect 55356 80332 55412 80388
rect 55244 79772 55300 79828
rect 56028 80556 56084 80612
rect 56364 80498 56420 80500
rect 56364 80446 56366 80498
rect 56366 80446 56418 80498
rect 56418 80446 56420 80498
rect 56364 80444 56420 80446
rect 56140 80220 56196 80276
rect 55916 79548 55972 79604
rect 54572 78988 54628 79044
rect 54236 78764 54292 78820
rect 52668 78034 52724 78036
rect 52668 77982 52670 78034
rect 52670 77982 52722 78034
rect 52722 77982 52724 78034
rect 52668 77980 52724 77982
rect 53116 77922 53172 77924
rect 53116 77870 53118 77922
rect 53118 77870 53170 77922
rect 53170 77870 53172 77922
rect 53116 77868 53172 77870
rect 52332 77196 52388 77252
rect 52892 77196 52948 77252
rect 52668 76188 52724 76244
rect 52668 75404 52724 75460
rect 52220 75068 52276 75124
rect 52892 74956 52948 75012
rect 52444 74172 52500 74228
rect 54236 77084 54292 77140
rect 53340 77026 53396 77028
rect 53340 76974 53342 77026
rect 53342 76974 53394 77026
rect 53394 76974 53396 77026
rect 53340 76972 53396 76974
rect 53788 77026 53844 77028
rect 53788 76974 53790 77026
rect 53790 76974 53842 77026
rect 53842 76974 53844 77026
rect 53788 76972 53844 76974
rect 54348 76972 54404 77028
rect 54236 76524 54292 76580
rect 53788 76300 53844 76356
rect 53564 76188 53620 76244
rect 53340 75180 53396 75236
rect 53676 74732 53732 74788
rect 53116 74172 53172 74228
rect 53340 74226 53396 74228
rect 53340 74174 53342 74226
rect 53342 74174 53394 74226
rect 53394 74174 53396 74226
rect 53340 74172 53396 74174
rect 54124 75122 54180 75124
rect 54124 75070 54126 75122
rect 54126 75070 54178 75122
rect 54178 75070 54180 75122
rect 54124 75068 54180 75070
rect 55244 76636 55300 76692
rect 54796 75180 54852 75236
rect 54908 76524 54964 76580
rect 54572 75068 54628 75124
rect 55132 75404 55188 75460
rect 55692 75122 55748 75124
rect 55692 75070 55694 75122
rect 55694 75070 55746 75122
rect 55746 75070 55748 75122
rect 55692 75068 55748 75070
rect 54348 75010 54404 75012
rect 54348 74958 54350 75010
rect 54350 74958 54402 75010
rect 54402 74958 54404 75010
rect 54348 74956 54404 74958
rect 54124 74844 54180 74900
rect 54460 74732 54516 74788
rect 54796 74732 54852 74788
rect 56588 81676 56644 81732
rect 57260 85202 57316 85204
rect 57260 85150 57262 85202
rect 57262 85150 57314 85202
rect 57314 85150 57316 85202
rect 57260 85148 57316 85150
rect 56924 84252 56980 84308
rect 57372 84194 57428 84196
rect 57372 84142 57374 84194
rect 57374 84142 57426 84194
rect 57426 84142 57428 84194
rect 57372 84140 57428 84142
rect 56924 82684 56980 82740
rect 57708 86044 57764 86100
rect 56924 80556 56980 80612
rect 56812 80386 56868 80388
rect 56812 80334 56814 80386
rect 56814 80334 56866 80386
rect 56866 80334 56868 80386
rect 56812 80332 56868 80334
rect 56700 79826 56756 79828
rect 56700 79774 56702 79826
rect 56702 79774 56754 79826
rect 56754 79774 56756 79826
rect 56700 79772 56756 79774
rect 56588 79548 56644 79604
rect 57036 80444 57092 80500
rect 57148 80386 57204 80388
rect 57148 80334 57150 80386
rect 57150 80334 57202 80386
rect 57202 80334 57204 80386
rect 57148 80332 57204 80334
rect 57372 80332 57428 80388
rect 57484 80444 57540 80500
rect 56924 79324 56980 79380
rect 57372 79660 57428 79716
rect 57596 80386 57652 80388
rect 57596 80334 57598 80386
rect 57598 80334 57650 80386
rect 57650 80334 57652 80386
rect 57596 80332 57652 80334
rect 58380 87218 58436 87220
rect 58380 87166 58382 87218
rect 58382 87166 58434 87218
rect 58434 87166 58436 87218
rect 58380 87164 58436 87166
rect 58716 86268 58772 86324
rect 58268 85986 58324 85988
rect 58268 85934 58270 85986
rect 58270 85934 58322 85986
rect 58322 85934 58324 85986
rect 58268 85932 58324 85934
rect 59948 86716 60004 86772
rect 59276 86268 59332 86324
rect 59836 85932 59892 85988
rect 59388 85314 59444 85316
rect 59388 85262 59390 85314
rect 59390 85262 59442 85314
rect 59442 85262 59444 85314
rect 59388 85260 59444 85262
rect 59500 85148 59556 85204
rect 58828 84306 58884 84308
rect 58828 84254 58830 84306
rect 58830 84254 58882 84306
rect 58882 84254 58884 84306
rect 58828 84252 58884 84254
rect 58940 82572 58996 82628
rect 58268 79602 58324 79604
rect 58268 79550 58270 79602
rect 58270 79550 58322 79602
rect 58322 79550 58324 79602
rect 58268 79548 58324 79550
rect 57932 79436 57988 79492
rect 57820 78540 57876 78596
rect 55916 74844 55972 74900
rect 55244 74732 55300 74788
rect 56476 76354 56532 76356
rect 56476 76302 56478 76354
rect 56478 76302 56530 76354
rect 56530 76302 56532 76354
rect 56476 76300 56532 76302
rect 56700 77868 56756 77924
rect 57372 77922 57428 77924
rect 57372 77870 57374 77922
rect 57374 77870 57426 77922
rect 57426 77870 57428 77922
rect 57372 77868 57428 77870
rect 57708 77250 57764 77252
rect 57708 77198 57710 77250
rect 57710 77198 57762 77250
rect 57762 77198 57764 77250
rect 57708 77196 57764 77198
rect 57372 76972 57428 77028
rect 57596 76578 57652 76580
rect 57596 76526 57598 76578
rect 57598 76526 57650 76578
rect 57650 76526 57652 76578
rect 57596 76524 57652 76526
rect 57372 76300 57428 76356
rect 58044 77980 58100 78036
rect 58156 77868 58212 77924
rect 58380 77644 58436 77700
rect 58156 76524 58212 76580
rect 58268 76636 58324 76692
rect 56476 74786 56532 74788
rect 56476 74734 56478 74786
rect 56478 74734 56530 74786
rect 56530 74734 56532 74786
rect 56476 74732 56532 74734
rect 51884 73218 51940 73220
rect 51884 73166 51886 73218
rect 51886 73166 51938 73218
rect 51938 73166 51940 73218
rect 51884 73164 51940 73166
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50428 71986 50484 71988
rect 50428 71934 50430 71986
rect 50430 71934 50482 71986
rect 50482 71934 50484 71986
rect 50428 71932 50484 71934
rect 50764 71538 50820 71540
rect 50764 71486 50766 71538
rect 50766 71486 50818 71538
rect 50818 71486 50820 71538
rect 50764 71484 50820 71486
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50204 68908 50260 68964
rect 49644 68572 49700 68628
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 50540 68402 50596 68404
rect 50540 68350 50542 68402
rect 50542 68350 50594 68402
rect 50594 68350 50596 68402
rect 50540 68348 50596 68350
rect 50988 68348 51044 68404
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 49756 67170 49812 67172
rect 49756 67118 49758 67170
rect 49758 67118 49810 67170
rect 49810 67118 49812 67170
rect 49756 67116 49812 67118
rect 48860 67058 48916 67060
rect 48860 67006 48862 67058
rect 48862 67006 48914 67058
rect 48914 67006 48916 67058
rect 48860 67004 48916 67006
rect 48300 66946 48356 66948
rect 48300 66894 48302 66946
rect 48302 66894 48354 66946
rect 48354 66894 48356 66946
rect 48300 66892 48356 66894
rect 49084 66892 49140 66948
rect 48860 63756 48916 63812
rect 48860 62188 48916 62244
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 47628 60508 47684 60564
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 46956 59218 47012 59220
rect 46956 59166 46958 59218
rect 46958 59166 47010 59218
rect 47010 59166 47012 59218
rect 46956 59164 47012 59166
rect 47964 59388 48020 59444
rect 47852 59330 47908 59332
rect 47852 59278 47854 59330
rect 47854 59278 47906 59330
rect 47906 59278 47908 59330
rect 47852 59276 47908 59278
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 2156 57036 2212 57092
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 47964 54236 48020 54292
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 48412 60898 48468 60900
rect 48412 60846 48414 60898
rect 48414 60846 48466 60898
rect 48466 60846 48468 60898
rect 48412 60844 48468 60846
rect 49308 66050 49364 66052
rect 49308 65998 49310 66050
rect 49310 65998 49362 66050
rect 49362 65998 49364 66050
rect 49308 65996 49364 65998
rect 49196 65660 49252 65716
rect 50428 67058 50484 67060
rect 50428 67006 50430 67058
rect 50430 67006 50482 67058
rect 50482 67006 50484 67058
rect 50428 67004 50484 67006
rect 50204 66892 50260 66948
rect 52332 73164 52388 73220
rect 53004 73164 53060 73220
rect 51436 71596 51492 71652
rect 52108 71650 52164 71652
rect 52108 71598 52110 71650
rect 52110 71598 52162 71650
rect 52162 71598 52164 71650
rect 52108 71596 52164 71598
rect 51212 68796 51268 68852
rect 52780 71596 52836 71652
rect 52556 71484 52612 71540
rect 52108 70476 52164 70532
rect 52668 70476 52724 70532
rect 51884 68626 51940 68628
rect 51884 68574 51886 68626
rect 51886 68574 51938 68626
rect 51938 68574 51940 68626
rect 51884 68572 51940 68574
rect 51100 67564 51156 67620
rect 52108 67564 52164 67620
rect 51100 67170 51156 67172
rect 51100 67118 51102 67170
rect 51102 67118 51154 67170
rect 51154 67118 51156 67170
rect 51100 67116 51156 67118
rect 50204 66162 50260 66164
rect 50204 66110 50206 66162
rect 50206 66110 50258 66162
rect 50258 66110 50260 66162
rect 50204 66108 50260 66110
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 50876 65660 50932 65716
rect 50540 65548 50596 65604
rect 49532 63756 49588 63812
rect 50988 64652 51044 64708
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 50316 63420 50372 63476
rect 49420 62860 49476 62916
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 50316 62188 50372 62244
rect 49420 60844 49476 60900
rect 51884 67170 51940 67172
rect 51884 67118 51886 67170
rect 51886 67118 51938 67170
rect 51938 67118 51940 67170
rect 51884 67116 51940 67118
rect 51660 66162 51716 66164
rect 51660 66110 51662 66162
rect 51662 66110 51714 66162
rect 51714 66110 51716 66162
rect 51660 66108 51716 66110
rect 51436 65548 51492 65604
rect 51772 65772 51828 65828
rect 52668 69356 52724 69412
rect 52668 69132 52724 69188
rect 52892 70194 52948 70196
rect 52892 70142 52894 70194
rect 52894 70142 52946 70194
rect 52946 70142 52948 70194
rect 52892 70140 52948 70142
rect 52780 68796 52836 68852
rect 53900 72492 53956 72548
rect 53340 70700 53396 70756
rect 53564 70700 53620 70756
rect 55468 72434 55524 72436
rect 55468 72382 55470 72434
rect 55470 72382 55522 72434
rect 55522 72382 55524 72434
rect 55468 72380 55524 72382
rect 54684 72322 54740 72324
rect 54684 72270 54686 72322
rect 54686 72270 54738 72322
rect 54738 72270 54740 72322
rect 54684 72268 54740 72270
rect 55244 72268 55300 72324
rect 53676 70476 53732 70532
rect 55132 70476 55188 70532
rect 54572 69916 54628 69972
rect 53676 69132 53732 69188
rect 52220 66050 52276 66052
rect 52220 65998 52222 66050
rect 52222 65998 52274 66050
rect 52274 65998 52276 66050
rect 52220 65996 52276 65998
rect 52556 66274 52612 66276
rect 52556 66222 52558 66274
rect 52558 66222 52610 66274
rect 52610 66222 52612 66274
rect 52556 66220 52612 66222
rect 52332 65884 52388 65940
rect 52108 65772 52164 65828
rect 52444 65772 52500 65828
rect 52444 65548 52500 65604
rect 52444 64594 52500 64596
rect 52444 64542 52446 64594
rect 52446 64542 52498 64594
rect 52498 64542 52500 64594
rect 52444 64540 52500 64542
rect 49756 60562 49812 60564
rect 49756 60510 49758 60562
rect 49758 60510 49810 60562
rect 49810 60510 49812 60562
rect 49756 60508 49812 60510
rect 48412 60002 48468 60004
rect 48412 59950 48414 60002
rect 48414 59950 48466 60002
rect 48466 59950 48468 60002
rect 48412 59948 48468 59950
rect 48748 59442 48804 59444
rect 48748 59390 48750 59442
rect 48750 59390 48802 59442
rect 48802 59390 48804 59442
rect 48748 59388 48804 59390
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50428 60732 50484 60788
rect 50764 60786 50820 60788
rect 50764 60734 50766 60786
rect 50766 60734 50818 60786
rect 50818 60734 50820 60786
rect 50764 60732 50820 60734
rect 51100 60732 51156 60788
rect 50876 60620 50932 60676
rect 50092 60060 50148 60116
rect 51212 60114 51268 60116
rect 51212 60062 51214 60114
rect 51214 60062 51266 60114
rect 51266 60062 51268 60114
rect 51212 60060 51268 60062
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 49196 59388 49252 59444
rect 50428 59388 50484 59444
rect 50316 59330 50372 59332
rect 50316 59278 50318 59330
rect 50318 59278 50370 59330
rect 50370 59278 50372 59330
rect 50316 59276 50372 59278
rect 48524 59218 48580 59220
rect 48524 59166 48526 59218
rect 48526 59166 48578 59218
rect 48578 59166 48580 59218
rect 48524 59164 48580 59166
rect 48524 58434 48580 58436
rect 48524 58382 48526 58434
rect 48526 58382 48578 58434
rect 48578 58382 48580 58434
rect 48524 58380 48580 58382
rect 49420 58434 49476 58436
rect 49420 58382 49422 58434
rect 49422 58382 49474 58434
rect 49474 58382 49476 58434
rect 49420 58380 49476 58382
rect 48300 56364 48356 56420
rect 48412 56252 48468 56308
rect 50540 58492 50596 58548
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50764 57484 50820 57540
rect 49756 56924 49812 56980
rect 49644 56364 49700 56420
rect 49532 56252 49588 56308
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50652 56306 50708 56308
rect 50652 56254 50654 56306
rect 50654 56254 50706 56306
rect 50706 56254 50708 56306
rect 50652 56252 50708 56254
rect 50204 55356 50260 55412
rect 51436 60674 51492 60676
rect 51436 60622 51438 60674
rect 51438 60622 51490 60674
rect 51490 60622 51492 60674
rect 51436 60620 51492 60622
rect 52444 63868 52500 63924
rect 52892 67564 52948 67620
rect 52892 67004 52948 67060
rect 52892 66220 52948 66276
rect 52780 63420 52836 63476
rect 53116 68348 53172 68404
rect 53340 67618 53396 67620
rect 53340 67566 53342 67618
rect 53342 67566 53394 67618
rect 53394 67566 53396 67618
rect 53340 67564 53396 67566
rect 53228 67116 53284 67172
rect 53116 65602 53172 65604
rect 53116 65550 53118 65602
rect 53118 65550 53170 65602
rect 53170 65550 53172 65602
rect 53116 65548 53172 65550
rect 53340 65660 53396 65716
rect 53676 68850 53732 68852
rect 53676 68798 53678 68850
rect 53678 68798 53730 68850
rect 53730 68798 53732 68850
rect 53676 68796 53732 68798
rect 56364 72716 56420 72772
rect 57820 73948 57876 74004
rect 56476 73164 56532 73220
rect 56140 72434 56196 72436
rect 56140 72382 56142 72434
rect 56142 72382 56194 72434
rect 56194 72382 56196 72434
rect 56140 72380 56196 72382
rect 57148 73836 57204 73892
rect 56476 72268 56532 72324
rect 56700 71650 56756 71652
rect 56700 71598 56702 71650
rect 56702 71598 56754 71650
rect 56754 71598 56756 71650
rect 56700 71596 56756 71598
rect 57260 71596 57316 71652
rect 58828 78876 58884 78932
rect 60508 87276 60564 87332
rect 60844 86940 60900 86996
rect 60508 85708 60564 85764
rect 60620 86770 60676 86772
rect 60620 86718 60622 86770
rect 60622 86718 60674 86770
rect 60674 86718 60676 86770
rect 60620 86716 60676 86718
rect 60396 85260 60452 85316
rect 60396 82626 60452 82628
rect 60396 82574 60398 82626
rect 60398 82574 60450 82626
rect 60450 82574 60452 82626
rect 60396 82572 60452 82574
rect 59724 81676 59780 81732
rect 60284 81730 60340 81732
rect 60284 81678 60286 81730
rect 60286 81678 60338 81730
rect 60338 81678 60340 81730
rect 60284 81676 60340 81678
rect 59500 79772 59556 79828
rect 62524 87836 62580 87892
rect 61852 87276 61908 87332
rect 62748 87500 62804 87556
rect 62412 87164 62468 87220
rect 62188 86770 62244 86772
rect 62188 86718 62190 86770
rect 62190 86718 62242 86770
rect 62242 86718 62244 86770
rect 62188 86716 62244 86718
rect 61516 86156 61572 86212
rect 60956 85762 61012 85764
rect 60956 85710 60958 85762
rect 60958 85710 61010 85762
rect 61010 85710 61012 85762
rect 60956 85708 61012 85710
rect 60844 82012 60900 82068
rect 59052 78988 59108 79044
rect 59500 79324 59556 79380
rect 58828 78316 58884 78372
rect 61740 85820 61796 85876
rect 63084 87164 63140 87220
rect 65916 88618 65972 88620
rect 65916 88566 65918 88618
rect 65918 88566 65970 88618
rect 65970 88566 65972 88618
rect 65916 88564 65972 88566
rect 66020 88618 66076 88620
rect 66020 88566 66022 88618
rect 66022 88566 66074 88618
rect 66074 88566 66076 88618
rect 66020 88564 66076 88566
rect 66124 88618 66180 88620
rect 66124 88566 66126 88618
rect 66126 88566 66178 88618
rect 66178 88566 66180 88618
rect 66124 88564 66180 88566
rect 63308 86716 63364 86772
rect 62412 85708 62468 85764
rect 62188 81900 62244 81956
rect 61516 80556 61572 80612
rect 61404 80498 61460 80500
rect 61404 80446 61406 80498
rect 61406 80446 61458 80498
rect 61458 80446 61460 80498
rect 61404 80444 61460 80446
rect 61180 79490 61236 79492
rect 61180 79438 61182 79490
rect 61182 79438 61234 79490
rect 61234 79438 61236 79490
rect 61180 79436 61236 79438
rect 60396 78818 60452 78820
rect 60396 78766 60398 78818
rect 60398 78766 60450 78818
rect 60450 78766 60452 78818
rect 60396 78764 60452 78766
rect 59724 78540 59780 78596
rect 60060 78034 60116 78036
rect 60060 77982 60062 78034
rect 60062 77982 60114 78034
rect 60114 77982 60116 78034
rect 60060 77980 60116 77982
rect 58604 77922 58660 77924
rect 58604 77870 58606 77922
rect 58606 77870 58658 77922
rect 58658 77870 58660 77922
rect 58604 77868 58660 77870
rect 58604 77026 58660 77028
rect 58604 76974 58606 77026
rect 58606 76974 58658 77026
rect 58658 76974 58660 77026
rect 58604 76972 58660 76974
rect 58940 76972 58996 77028
rect 58492 76466 58548 76468
rect 58492 76414 58494 76466
rect 58494 76414 58546 76466
rect 58546 76414 58548 76466
rect 58492 76412 58548 76414
rect 58156 73948 58212 74004
rect 58940 76412 58996 76468
rect 58268 73836 58324 73892
rect 59724 74002 59780 74004
rect 59724 73950 59726 74002
rect 59726 73950 59778 74002
rect 59778 73950 59780 74002
rect 59724 73948 59780 73950
rect 60396 74114 60452 74116
rect 60396 74062 60398 74114
rect 60398 74062 60450 74114
rect 60450 74062 60452 74114
rect 60396 74060 60452 74062
rect 58044 72770 58100 72772
rect 58044 72718 58046 72770
rect 58046 72718 58098 72770
rect 58098 72718 58100 72770
rect 58044 72716 58100 72718
rect 57820 72492 57876 72548
rect 58380 72546 58436 72548
rect 58380 72494 58382 72546
rect 58382 72494 58434 72546
rect 58434 72494 58436 72546
rect 58380 72492 58436 72494
rect 59500 73836 59556 73892
rect 57932 71090 57988 71092
rect 57932 71038 57934 71090
rect 57934 71038 57986 71090
rect 57986 71038 57988 71090
rect 57932 71036 57988 71038
rect 57372 70588 57428 70644
rect 56476 70476 56532 70532
rect 56252 70364 56308 70420
rect 55580 70140 55636 70196
rect 54684 68684 54740 68740
rect 53788 67618 53844 67620
rect 53788 67566 53790 67618
rect 53790 67566 53842 67618
rect 53842 67566 53844 67618
rect 53788 67564 53844 67566
rect 54236 67452 54292 67508
rect 53788 67170 53844 67172
rect 53788 67118 53790 67170
rect 53790 67118 53842 67170
rect 53842 67118 53844 67170
rect 53788 67116 53844 67118
rect 54684 66780 54740 66836
rect 54012 65884 54068 65940
rect 54124 65602 54180 65604
rect 54124 65550 54126 65602
rect 54126 65550 54178 65602
rect 54178 65550 54180 65602
rect 54124 65548 54180 65550
rect 54572 65490 54628 65492
rect 54572 65438 54574 65490
rect 54574 65438 54626 65490
rect 54626 65438 54628 65490
rect 54572 65436 54628 65438
rect 53452 64876 53508 64932
rect 53340 64706 53396 64708
rect 53340 64654 53342 64706
rect 53342 64654 53394 64706
rect 53394 64654 53396 64706
rect 53340 64652 53396 64654
rect 53676 65212 53732 65268
rect 54124 64876 54180 64932
rect 53676 64540 53732 64596
rect 54684 64540 54740 64596
rect 53004 63420 53060 63476
rect 52220 63084 52276 63140
rect 52668 63250 52724 63252
rect 52668 63198 52670 63250
rect 52670 63198 52722 63250
rect 52722 63198 52724 63250
rect 52668 63196 52724 63198
rect 51772 62860 51828 62916
rect 51772 62412 51828 62468
rect 53340 63196 53396 63252
rect 53452 63810 53508 63812
rect 53452 63758 53454 63810
rect 53454 63758 53506 63810
rect 53506 63758 53508 63810
rect 53452 63756 53508 63758
rect 52668 62466 52724 62468
rect 52668 62414 52670 62466
rect 52670 62414 52722 62466
rect 52722 62414 52724 62466
rect 52668 62412 52724 62414
rect 53564 63084 53620 63140
rect 54236 63922 54292 63924
rect 54236 63870 54238 63922
rect 54238 63870 54290 63922
rect 54290 63870 54292 63922
rect 54236 63868 54292 63870
rect 54460 63308 54516 63364
rect 52332 61292 52388 61348
rect 51884 60732 51940 60788
rect 51772 60002 51828 60004
rect 51772 59950 51774 60002
rect 51774 59950 51826 60002
rect 51826 59950 51828 60002
rect 51772 59948 51828 59950
rect 51996 58546 52052 58548
rect 51996 58494 51998 58546
rect 51998 58494 52050 58546
rect 52050 58494 52052 58546
rect 51996 58492 52052 58494
rect 51212 56978 51268 56980
rect 51212 56926 51214 56978
rect 51214 56926 51266 56978
rect 51266 56926 51268 56978
rect 51212 56924 51268 56926
rect 51996 56924 52052 56980
rect 51436 56252 51492 56308
rect 51212 55410 51268 55412
rect 51212 55358 51214 55410
rect 51214 55358 51266 55410
rect 51266 55358 51268 55410
rect 51212 55356 51268 55358
rect 52220 57538 52276 57540
rect 52220 57486 52222 57538
rect 52222 57486 52274 57538
rect 52274 57486 52276 57538
rect 52220 57484 52276 57486
rect 52108 55186 52164 55188
rect 52108 55134 52110 55186
rect 52110 55134 52162 55186
rect 52162 55134 52164 55186
rect 52108 55132 52164 55134
rect 52220 56252 52276 56308
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 48188 53618 48244 53620
rect 48188 53566 48190 53618
rect 48190 53566 48242 53618
rect 48242 53566 48244 53618
rect 48188 53564 48244 53566
rect 48860 52892 48916 52948
rect 49532 53618 49588 53620
rect 49532 53566 49534 53618
rect 49534 53566 49586 53618
rect 49586 53566 49588 53618
rect 49532 53564 49588 53566
rect 50988 54514 51044 54516
rect 50988 54462 50990 54514
rect 50990 54462 51042 54514
rect 51042 54462 51044 54514
rect 50988 54460 51044 54462
rect 51772 54290 51828 54292
rect 51772 54238 51774 54290
rect 51774 54238 51826 54290
rect 51826 54238 51828 54290
rect 51772 54236 51828 54238
rect 51660 53676 51716 53732
rect 52444 60620 52500 60676
rect 52780 60002 52836 60004
rect 52780 59950 52782 60002
rect 52782 59950 52834 60002
rect 52834 59950 52836 60002
rect 52780 59948 52836 59950
rect 52444 58940 52500 58996
rect 53004 57650 53060 57652
rect 53004 57598 53006 57650
rect 53006 57598 53058 57650
rect 53058 57598 53060 57650
rect 53004 57596 53060 57598
rect 52668 56252 52724 56308
rect 52780 57484 52836 57540
rect 50876 53452 50932 53508
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 52108 53116 52164 53172
rect 52444 55132 52500 55188
rect 49532 52946 49588 52948
rect 49532 52894 49534 52946
rect 49534 52894 49586 52946
rect 49586 52894 49588 52946
rect 49532 52892 49588 52894
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50988 50540 51044 50596
rect 48076 49980 48132 50036
rect 50428 50428 50484 50484
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 49868 49420 49924 49476
rect 51548 50594 51604 50596
rect 51548 50542 51550 50594
rect 51550 50542 51602 50594
rect 51602 50542 51604 50594
rect 51548 50540 51604 50542
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 50428 48748 50484 48804
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 50092 47570 50148 47572
rect 50092 47518 50094 47570
rect 50094 47518 50146 47570
rect 50146 47518 50148 47570
rect 50092 47516 50148 47518
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 48748 44156 48804 44212
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 49756 44210 49812 44212
rect 49756 44158 49758 44210
rect 49758 44158 49810 44210
rect 49810 44158 49812 44210
rect 49756 44156 49812 44158
rect 49084 44044 49140 44100
rect 50092 44044 50148 44100
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 51884 50370 51940 50372
rect 51884 50318 51886 50370
rect 51886 50318 51938 50370
rect 51938 50318 51940 50370
rect 51884 50316 51940 50318
rect 51884 49420 51940 49476
rect 53116 55468 53172 55524
rect 52780 54514 52836 54516
rect 52780 54462 52782 54514
rect 52782 54462 52834 54514
rect 52834 54462 52836 54514
rect 52780 54460 52836 54462
rect 52780 54012 52836 54068
rect 53004 53676 53060 53732
rect 52556 53506 52612 53508
rect 52556 53454 52558 53506
rect 52558 53454 52610 53506
rect 52610 53454 52612 53506
rect 52556 53452 52612 53454
rect 52892 53170 52948 53172
rect 52892 53118 52894 53170
rect 52894 53118 52946 53170
rect 52946 53118 52948 53170
rect 52892 53116 52948 53118
rect 53004 52892 53060 52948
rect 53116 54460 53172 54516
rect 52556 52108 52612 52164
rect 52892 52220 52948 52276
rect 52332 50652 52388 50708
rect 52332 50482 52388 50484
rect 52332 50430 52334 50482
rect 52334 50430 52386 50482
rect 52386 50430 52388 50482
rect 52332 50428 52388 50430
rect 48524 43538 48580 43540
rect 48524 43486 48526 43538
rect 48526 43486 48578 43538
rect 48578 43486 48580 43538
rect 48524 43484 48580 43486
rect 49756 43538 49812 43540
rect 49756 43486 49758 43538
rect 49758 43486 49810 43538
rect 49810 43486 49812 43538
rect 49756 43484 49812 43486
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 50092 43426 50148 43428
rect 50092 43374 50094 43426
rect 50094 43374 50146 43426
rect 50146 43374 50148 43426
rect 50092 43372 50148 43374
rect 50876 43538 50932 43540
rect 50876 43486 50878 43538
rect 50878 43486 50930 43538
rect 50930 43486 50932 43538
rect 50876 43484 50932 43486
rect 50764 43260 50820 43316
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 49532 41074 49588 41076
rect 49532 41022 49534 41074
rect 49534 41022 49586 41074
rect 49586 41022 49588 41074
rect 49532 41020 49588 41022
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 14252 39340 14308 39396
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 1820 37490 1876 37492
rect 1820 37438 1822 37490
rect 1822 37438 1874 37490
rect 1874 37438 1876 37490
rect 1820 37436 1876 37438
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2156 12738 2212 12740
rect 2156 12686 2158 12738
rect 2158 12686 2210 12738
rect 2210 12686 2212 12738
rect 2156 12684 2212 12686
rect 1820 12460 1876 12516
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 6972 3330 7028 3332
rect 6972 3278 6974 3330
rect 6974 3278 7026 3330
rect 7026 3278 7028 3330
rect 6972 3276 7028 3278
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50764 41186 50820 41188
rect 50764 41134 50766 41186
rect 50766 41134 50818 41186
rect 50818 41134 50820 41186
rect 50764 41132 50820 41134
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 51996 43426 52052 43428
rect 51996 43374 51998 43426
rect 51998 43374 52050 43426
rect 52050 43374 52052 43426
rect 51996 43372 52052 43374
rect 51772 41804 51828 41860
rect 51436 41074 51492 41076
rect 51436 41022 51438 41074
rect 51438 41022 51490 41074
rect 51490 41022 51492 41074
rect 51436 41020 51492 41022
rect 50540 39394 50596 39396
rect 50540 39342 50542 39394
rect 50542 39342 50594 39394
rect 50594 39342 50596 39394
rect 50540 39340 50596 39342
rect 51436 39506 51492 39508
rect 51436 39454 51438 39506
rect 51438 39454 51490 39506
rect 51490 39454 51492 39506
rect 51436 39452 51492 39454
rect 51100 39340 51156 39396
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 52668 49868 52724 49924
rect 52444 48412 52500 48468
rect 52556 49420 52612 49476
rect 52220 48300 52276 48356
rect 52668 49138 52724 49140
rect 52668 49086 52670 49138
rect 52670 49086 52722 49138
rect 52722 49086 52724 49138
rect 52668 49084 52724 49086
rect 52780 48524 52836 48580
rect 52668 48130 52724 48132
rect 52668 48078 52670 48130
rect 52670 48078 52722 48130
rect 52722 48078 52724 48130
rect 52668 48076 52724 48078
rect 54460 63138 54516 63140
rect 54460 63086 54462 63138
rect 54462 63086 54514 63138
rect 54514 63086 54516 63138
rect 54460 63084 54516 63086
rect 54124 62636 54180 62692
rect 53340 61346 53396 61348
rect 53340 61294 53342 61346
rect 53342 61294 53394 61346
rect 53394 61294 53396 61346
rect 53340 61292 53396 61294
rect 55244 66332 55300 66388
rect 55020 65602 55076 65604
rect 55020 65550 55022 65602
rect 55022 65550 55074 65602
rect 55074 65550 55076 65602
rect 55020 65548 55076 65550
rect 55356 65490 55412 65492
rect 55356 65438 55358 65490
rect 55358 65438 55410 65490
rect 55410 65438 55412 65490
rect 55356 65436 55412 65438
rect 55356 64316 55412 64372
rect 55020 63868 55076 63924
rect 55132 62524 55188 62580
rect 55692 69468 55748 69524
rect 56476 69522 56532 69524
rect 56476 69470 56478 69522
rect 56478 69470 56530 69522
rect 56530 69470 56532 69522
rect 56476 69468 56532 69470
rect 57148 69468 57204 69524
rect 56476 69244 56532 69300
rect 57596 69970 57652 69972
rect 57596 69918 57598 69970
rect 57598 69918 57650 69970
rect 57650 69918 57652 69970
rect 57596 69916 57652 69918
rect 57932 69580 57988 69636
rect 57820 69298 57876 69300
rect 57820 69246 57822 69298
rect 57822 69246 57874 69298
rect 57874 69246 57876 69298
rect 57820 69244 57876 69246
rect 56476 66386 56532 66388
rect 56476 66334 56478 66386
rect 56478 66334 56530 66386
rect 56530 66334 56532 66386
rect 56476 66332 56532 66334
rect 58044 66332 58100 66388
rect 55804 66220 55860 66276
rect 55804 65490 55860 65492
rect 55804 65438 55806 65490
rect 55806 65438 55858 65490
rect 55858 65438 55860 65490
rect 55804 65436 55860 65438
rect 56364 64818 56420 64820
rect 56364 64766 56366 64818
rect 56366 64766 56418 64818
rect 56418 64766 56420 64818
rect 56364 64764 56420 64766
rect 55692 63420 55748 63476
rect 56476 64482 56532 64484
rect 56476 64430 56478 64482
rect 56478 64430 56530 64482
rect 56530 64430 56532 64482
rect 56476 64428 56532 64430
rect 56924 64204 56980 64260
rect 56364 63420 56420 63476
rect 56140 61516 56196 61572
rect 55020 61458 55076 61460
rect 55020 61406 55022 61458
rect 55022 61406 55074 61458
rect 55074 61406 55076 61458
rect 55020 61404 55076 61406
rect 55692 61458 55748 61460
rect 55692 61406 55694 61458
rect 55694 61406 55746 61458
rect 55746 61406 55748 61458
rect 55692 61404 55748 61406
rect 55132 61346 55188 61348
rect 55132 61294 55134 61346
rect 55134 61294 55186 61346
rect 55186 61294 55188 61346
rect 55132 61292 55188 61294
rect 56140 61346 56196 61348
rect 56140 61294 56142 61346
rect 56142 61294 56194 61346
rect 56194 61294 56196 61346
rect 56140 61292 56196 61294
rect 56700 62636 56756 62692
rect 53676 60002 53732 60004
rect 53676 59950 53678 60002
rect 53678 59950 53730 60002
rect 53730 59950 53732 60002
rect 53676 59948 53732 59950
rect 53340 56924 53396 56980
rect 53564 56252 53620 56308
rect 54236 59164 54292 59220
rect 54348 59612 54404 59668
rect 54460 59388 54516 59444
rect 56140 60786 56196 60788
rect 56140 60734 56142 60786
rect 56142 60734 56194 60786
rect 56194 60734 56196 60786
rect 56140 60732 56196 60734
rect 55580 60172 55636 60228
rect 56924 63084 56980 63140
rect 57596 64652 57652 64708
rect 57484 64594 57540 64596
rect 57484 64542 57486 64594
rect 57486 64542 57538 64594
rect 57538 64542 57540 64594
rect 57484 64540 57540 64542
rect 57820 64594 57876 64596
rect 57820 64542 57822 64594
rect 57822 64542 57874 64594
rect 57874 64542 57876 64594
rect 57820 64540 57876 64542
rect 57596 64316 57652 64372
rect 57484 64034 57540 64036
rect 57484 63982 57486 64034
rect 57486 63982 57538 64034
rect 57538 63982 57540 64034
rect 57484 63980 57540 63982
rect 57036 62636 57092 62692
rect 57372 63308 57428 63364
rect 57596 63420 57652 63476
rect 57708 63308 57764 63364
rect 58492 71596 58548 71652
rect 58604 70364 58660 70420
rect 59052 71036 59108 71092
rect 58828 70140 58884 70196
rect 58716 70028 58772 70084
rect 59500 71036 59556 71092
rect 60396 72546 60452 72548
rect 60396 72494 60398 72546
rect 60398 72494 60450 72546
rect 60450 72494 60452 72546
rect 60396 72492 60452 72494
rect 60284 70588 60340 70644
rect 61292 78594 61348 78596
rect 61292 78542 61294 78594
rect 61294 78542 61346 78594
rect 61346 78542 61348 78594
rect 61292 78540 61348 78542
rect 60956 78316 61012 78372
rect 61740 78316 61796 78372
rect 63420 86156 63476 86212
rect 63084 85874 63140 85876
rect 63084 85822 63086 85874
rect 63086 85822 63138 85874
rect 63138 85822 63140 85874
rect 63084 85820 63140 85822
rect 62972 85708 63028 85764
rect 63756 87218 63812 87220
rect 63756 87166 63758 87218
rect 63758 87166 63810 87218
rect 63810 87166 63812 87218
rect 63756 87164 63812 87166
rect 64428 87836 64484 87892
rect 64316 87554 64372 87556
rect 64316 87502 64318 87554
rect 64318 87502 64370 87554
rect 64370 87502 64372 87554
rect 64316 87500 64372 87502
rect 64540 86268 64596 86324
rect 63868 85708 63924 85764
rect 64316 85762 64372 85764
rect 64316 85710 64318 85762
rect 64318 85710 64370 85762
rect 64370 85710 64372 85762
rect 64316 85708 64372 85710
rect 63756 84812 63812 84868
rect 64316 84306 64372 84308
rect 64316 84254 64318 84306
rect 64318 84254 64370 84306
rect 64370 84254 64372 84306
rect 64316 84252 64372 84254
rect 64428 84028 64484 84084
rect 62524 81900 62580 81956
rect 62636 80556 62692 80612
rect 67452 87276 67508 87332
rect 65916 87050 65972 87052
rect 65916 86998 65918 87050
rect 65918 86998 65970 87050
rect 65970 86998 65972 87050
rect 65916 86996 65972 86998
rect 66020 87050 66076 87052
rect 66020 86998 66022 87050
rect 66022 86998 66074 87050
rect 66074 86998 66076 87050
rect 66020 86996 66076 86998
rect 66124 87050 66180 87052
rect 66124 86998 66126 87050
rect 66126 86998 66178 87050
rect 66178 86998 66180 87050
rect 66124 86996 66180 86998
rect 65548 86380 65604 86436
rect 65772 86268 65828 86324
rect 65772 85820 65828 85876
rect 66668 86434 66724 86436
rect 66668 86382 66670 86434
rect 66670 86382 66722 86434
rect 66722 86382 66724 86434
rect 66668 86380 66724 86382
rect 65436 85762 65492 85764
rect 65436 85710 65438 85762
rect 65438 85710 65490 85762
rect 65490 85710 65492 85762
rect 65436 85708 65492 85710
rect 65916 85482 65972 85484
rect 65916 85430 65918 85482
rect 65918 85430 65970 85482
rect 65970 85430 65972 85482
rect 65916 85428 65972 85430
rect 66020 85482 66076 85484
rect 66020 85430 66022 85482
rect 66022 85430 66074 85482
rect 66074 85430 66076 85482
rect 66020 85428 66076 85430
rect 66124 85482 66180 85484
rect 66124 85430 66126 85482
rect 66126 85430 66178 85482
rect 66178 85430 66180 85482
rect 66124 85428 66180 85430
rect 65100 84028 65156 84084
rect 65772 84530 65828 84532
rect 65772 84478 65774 84530
rect 65774 84478 65826 84530
rect 65826 84478 65828 84530
rect 65772 84476 65828 84478
rect 63980 82066 64036 82068
rect 63980 82014 63982 82066
rect 63982 82014 64034 82066
rect 64034 82014 64036 82066
rect 63980 82012 64036 82014
rect 63644 81900 63700 81956
rect 62972 80444 63028 80500
rect 63420 81676 63476 81732
rect 64092 81676 64148 81732
rect 63420 80556 63476 80612
rect 63644 80668 63700 80724
rect 64428 81730 64484 81732
rect 64428 81678 64430 81730
rect 64430 81678 64482 81730
rect 64482 81678 64484 81730
rect 64428 81676 64484 81678
rect 64204 80668 64260 80724
rect 62636 79548 62692 79604
rect 62300 78818 62356 78820
rect 62300 78766 62302 78818
rect 62302 78766 62354 78818
rect 62354 78766 62356 78818
rect 62300 78764 62356 78766
rect 63308 79602 63364 79604
rect 63308 79550 63310 79602
rect 63310 79550 63362 79602
rect 63362 79550 63364 79602
rect 63308 79548 63364 79550
rect 61628 77644 61684 77700
rect 61516 75852 61572 75908
rect 60620 74898 60676 74900
rect 60620 74846 60622 74898
rect 60622 74846 60674 74898
rect 60674 74846 60676 74898
rect 60620 74844 60676 74846
rect 61516 74732 61572 74788
rect 61516 74114 61572 74116
rect 61516 74062 61518 74114
rect 61518 74062 61570 74114
rect 61570 74062 61572 74114
rect 61516 74060 61572 74062
rect 61516 73500 61572 73556
rect 60844 73218 60900 73220
rect 60844 73166 60846 73218
rect 60846 73166 60898 73218
rect 60898 73166 60900 73218
rect 60844 73164 60900 73166
rect 60620 71036 60676 71092
rect 60956 71148 61012 71204
rect 60620 70364 60676 70420
rect 59276 70194 59332 70196
rect 59276 70142 59278 70194
rect 59278 70142 59330 70194
rect 59330 70142 59332 70194
rect 59276 70140 59332 70142
rect 58716 68796 58772 68852
rect 59724 70082 59780 70084
rect 59724 70030 59726 70082
rect 59726 70030 59778 70082
rect 59778 70030 59780 70082
rect 59724 70028 59780 70030
rect 57932 64092 57988 64148
rect 58044 64706 58100 64708
rect 58044 64654 58046 64706
rect 58046 64654 58098 64706
rect 58098 64654 58100 64706
rect 58044 64652 58100 64654
rect 57932 63922 57988 63924
rect 57932 63870 57934 63922
rect 57934 63870 57986 63922
rect 57986 63870 57988 63922
rect 57932 63868 57988 63870
rect 58828 66162 58884 66164
rect 58828 66110 58830 66162
rect 58830 66110 58882 66162
rect 58882 66110 58884 66162
rect 58828 66108 58884 66110
rect 58828 65772 58884 65828
rect 59052 65772 59108 65828
rect 58940 65490 58996 65492
rect 58940 65438 58942 65490
rect 58942 65438 58994 65490
rect 58994 65438 58996 65490
rect 58940 65436 58996 65438
rect 58492 64316 58548 64372
rect 57820 62300 57876 62356
rect 58156 63308 58212 63364
rect 58268 63250 58324 63252
rect 58268 63198 58270 63250
rect 58270 63198 58322 63250
rect 58322 63198 58324 63250
rect 58268 63196 58324 63198
rect 59500 64652 59556 64708
rect 59612 65436 59668 65492
rect 59388 64594 59444 64596
rect 59388 64542 59390 64594
rect 59390 64542 59442 64594
rect 59442 64542 59444 64594
rect 59388 64540 59444 64542
rect 58716 63980 58772 64036
rect 58604 62524 58660 62580
rect 58604 62354 58660 62356
rect 58604 62302 58606 62354
rect 58606 62302 58658 62354
rect 58658 62302 58660 62354
rect 58604 62300 58660 62302
rect 56476 59500 56532 59556
rect 56812 59836 56868 59892
rect 57036 61292 57092 61348
rect 56812 59276 56868 59332
rect 55468 58828 55524 58884
rect 54460 58604 54516 58660
rect 55244 58434 55300 58436
rect 55244 58382 55246 58434
rect 55246 58382 55298 58434
rect 55298 58382 55300 58434
rect 55244 58380 55300 58382
rect 54684 58322 54740 58324
rect 54684 58270 54686 58322
rect 54686 58270 54738 58322
rect 54738 58270 54740 58322
rect 54684 58268 54740 58270
rect 55916 58322 55972 58324
rect 55916 58270 55918 58322
rect 55918 58270 55970 58322
rect 55970 58270 55972 58322
rect 55916 58268 55972 58270
rect 54348 56978 54404 56980
rect 54348 56926 54350 56978
rect 54350 56926 54402 56978
rect 54402 56926 54404 56978
rect 54348 56924 54404 56926
rect 54460 56364 54516 56420
rect 56700 57036 56756 57092
rect 56476 56700 56532 56756
rect 54572 56252 54628 56308
rect 56588 56588 56644 56644
rect 56476 56082 56532 56084
rect 56476 56030 56478 56082
rect 56478 56030 56530 56082
rect 56530 56030 56532 56082
rect 56476 56028 56532 56030
rect 55468 55468 55524 55524
rect 55020 54514 55076 54516
rect 55020 54462 55022 54514
rect 55022 54462 55074 54514
rect 55074 54462 55076 54514
rect 55020 54460 55076 54462
rect 53452 54012 53508 54068
rect 53900 54012 53956 54068
rect 55132 52892 55188 52948
rect 53340 52274 53396 52276
rect 53340 52222 53342 52274
rect 53342 52222 53394 52274
rect 53394 52222 53396 52274
rect 53340 52220 53396 52222
rect 54348 51884 54404 51940
rect 54124 51660 54180 51716
rect 53676 50652 53732 50708
rect 53004 50316 53060 50372
rect 53564 50370 53620 50372
rect 53564 50318 53566 50370
rect 53566 50318 53618 50370
rect 53618 50318 53620 50370
rect 53564 50316 53620 50318
rect 54348 50540 54404 50596
rect 55020 51884 55076 51940
rect 54908 50652 54964 50708
rect 54572 50370 54628 50372
rect 54572 50318 54574 50370
rect 54574 50318 54626 50370
rect 54626 50318 54628 50370
rect 54572 50316 54628 50318
rect 54348 49756 54404 49812
rect 54460 49532 54516 49588
rect 54124 49084 54180 49140
rect 53340 48802 53396 48804
rect 53340 48750 53342 48802
rect 53342 48750 53394 48802
rect 53394 48750 53396 48802
rect 53340 48748 53396 48750
rect 53564 48802 53620 48804
rect 53564 48750 53566 48802
rect 53566 48750 53618 48802
rect 53618 48750 53620 48802
rect 53564 48748 53620 48750
rect 53116 47516 53172 47572
rect 52892 45276 52948 45332
rect 53452 48412 53508 48468
rect 55580 55244 55636 55300
rect 59276 64316 59332 64372
rect 58940 63980 58996 64036
rect 59052 64092 59108 64148
rect 58940 63084 58996 63140
rect 59500 63532 59556 63588
rect 58828 62860 58884 62916
rect 59836 69468 59892 69524
rect 60732 70140 60788 70196
rect 60396 69522 60452 69524
rect 60396 69470 60398 69522
rect 60398 69470 60450 69522
rect 60450 69470 60452 69522
rect 60396 69468 60452 69470
rect 60732 68908 60788 68964
rect 60620 67730 60676 67732
rect 60620 67678 60622 67730
rect 60622 67678 60674 67730
rect 60674 67678 60676 67730
rect 60620 67676 60676 67678
rect 60396 66274 60452 66276
rect 60396 66222 60398 66274
rect 60398 66222 60450 66274
rect 60450 66222 60452 66274
rect 60396 66220 60452 66222
rect 60508 66108 60564 66164
rect 61516 70364 61572 70420
rect 60956 70028 61012 70084
rect 61516 68626 61572 68628
rect 61516 68574 61518 68626
rect 61518 68574 61570 68626
rect 61570 68574 61572 68626
rect 61516 68572 61572 68574
rect 61516 67730 61572 67732
rect 61516 67678 61518 67730
rect 61518 67678 61570 67730
rect 61570 67678 61572 67730
rect 61516 67676 61572 67678
rect 62076 77250 62132 77252
rect 62076 77198 62078 77250
rect 62078 77198 62130 77250
rect 62130 77198 62132 77250
rect 62076 77196 62132 77198
rect 62972 78540 63028 78596
rect 63420 78316 63476 78372
rect 63084 77308 63140 77364
rect 62972 77196 63028 77252
rect 63532 76690 63588 76692
rect 63532 76638 63534 76690
rect 63534 76638 63586 76690
rect 63586 76638 63588 76690
rect 63532 76636 63588 76638
rect 63868 76354 63924 76356
rect 63868 76302 63870 76354
rect 63870 76302 63922 76354
rect 63922 76302 63924 76354
rect 63868 76300 63924 76302
rect 66220 84866 66276 84868
rect 66220 84814 66222 84866
rect 66222 84814 66274 84866
rect 66274 84814 66276 84866
rect 66220 84812 66276 84814
rect 65916 83914 65972 83916
rect 65916 83862 65918 83914
rect 65918 83862 65970 83914
rect 65970 83862 65972 83914
rect 65916 83860 65972 83862
rect 66020 83914 66076 83916
rect 66020 83862 66022 83914
rect 66022 83862 66074 83914
rect 66074 83862 66076 83914
rect 66020 83860 66076 83862
rect 66124 83914 66180 83916
rect 66124 83862 66126 83914
rect 66126 83862 66178 83914
rect 66178 83862 66180 83914
rect 66124 83860 66180 83862
rect 65916 82346 65972 82348
rect 65916 82294 65918 82346
rect 65918 82294 65970 82346
rect 65970 82294 65972 82346
rect 65916 82292 65972 82294
rect 66020 82346 66076 82348
rect 66020 82294 66022 82346
rect 66022 82294 66074 82346
rect 66074 82294 66076 82346
rect 66020 82292 66076 82294
rect 66124 82346 66180 82348
rect 66124 82294 66126 82346
rect 66126 82294 66178 82346
rect 66178 82294 66180 82346
rect 66124 82292 66180 82294
rect 65772 81340 65828 81396
rect 67228 85820 67284 85876
rect 67116 84924 67172 84980
rect 68236 87276 68292 87332
rect 69244 86604 69300 86660
rect 68572 86546 68628 86548
rect 68572 86494 68574 86546
rect 68574 86494 68626 86546
rect 68626 86494 68628 86546
rect 68572 86492 68628 86494
rect 67452 85708 67508 85764
rect 68348 86380 68404 86436
rect 67340 84924 67396 84980
rect 66556 84476 66612 84532
rect 67116 84418 67172 84420
rect 67116 84366 67118 84418
rect 67118 84366 67170 84418
rect 67170 84366 67172 84418
rect 67116 84364 67172 84366
rect 66444 84252 66500 84308
rect 68012 84364 68068 84420
rect 67340 84028 67396 84084
rect 67676 84028 67732 84084
rect 68684 82236 68740 82292
rect 66332 81340 66388 81396
rect 65916 80778 65972 80780
rect 65916 80726 65918 80778
rect 65918 80726 65970 80778
rect 65970 80726 65972 80778
rect 65916 80724 65972 80726
rect 66020 80778 66076 80780
rect 66020 80726 66022 80778
rect 66022 80726 66074 80778
rect 66074 80726 66076 80778
rect 66020 80724 66076 80726
rect 66124 80778 66180 80780
rect 66124 80726 66126 80778
rect 66126 80726 66178 80778
rect 66178 80726 66180 80778
rect 66124 80724 66180 80726
rect 68012 80332 68068 80388
rect 68124 81004 68180 81060
rect 66444 79714 66500 79716
rect 66444 79662 66446 79714
rect 66446 79662 66498 79714
rect 66498 79662 66500 79714
rect 66444 79660 66500 79662
rect 65660 79548 65716 79604
rect 65916 79210 65972 79212
rect 65916 79158 65918 79210
rect 65918 79158 65970 79210
rect 65970 79158 65972 79210
rect 65916 79156 65972 79158
rect 66020 79210 66076 79212
rect 66020 79158 66022 79210
rect 66022 79158 66074 79210
rect 66074 79158 66076 79210
rect 66020 79156 66076 79158
rect 66124 79210 66180 79212
rect 66124 79158 66126 79210
rect 66126 79158 66178 79210
rect 66178 79158 66180 79210
rect 66124 79156 66180 79158
rect 66332 78876 66388 78932
rect 66780 79436 66836 79492
rect 66556 78764 66612 78820
rect 67228 78930 67284 78932
rect 67228 78878 67230 78930
rect 67230 78878 67282 78930
rect 67282 78878 67284 78930
rect 67228 78876 67284 78878
rect 62972 75794 63028 75796
rect 62972 75742 62974 75794
rect 62974 75742 63026 75794
rect 63026 75742 63028 75794
rect 62972 75740 63028 75742
rect 61852 73948 61908 74004
rect 62076 73164 62132 73220
rect 63868 75740 63924 75796
rect 62524 72940 62580 72996
rect 61740 72546 61796 72548
rect 61740 72494 61742 72546
rect 61742 72494 61794 72546
rect 61794 72494 61796 72546
rect 61740 72492 61796 72494
rect 62188 71090 62244 71092
rect 62188 71038 62190 71090
rect 62190 71038 62242 71090
rect 62242 71038 62244 71090
rect 62188 71036 62244 71038
rect 62188 68626 62244 68628
rect 62188 68574 62190 68626
rect 62190 68574 62242 68626
rect 62242 68574 62244 68626
rect 62188 68572 62244 68574
rect 62300 68460 62356 68516
rect 61852 68348 61908 68404
rect 60844 64988 60900 65044
rect 62748 72156 62804 72212
rect 62748 71596 62804 71652
rect 63644 72156 63700 72212
rect 65436 76972 65492 77028
rect 65916 77642 65972 77644
rect 65916 77590 65918 77642
rect 65918 77590 65970 77642
rect 65970 77590 65972 77642
rect 65916 77588 65972 77590
rect 66020 77642 66076 77644
rect 66020 77590 66022 77642
rect 66022 77590 66074 77642
rect 66074 77590 66076 77642
rect 66020 77588 66076 77590
rect 66124 77642 66180 77644
rect 66124 77590 66126 77642
rect 66126 77590 66178 77642
rect 66178 77590 66180 77642
rect 66124 77588 66180 77590
rect 64540 76690 64596 76692
rect 64540 76638 64542 76690
rect 64542 76638 64594 76690
rect 64594 76638 64596 76690
rect 64540 76636 64596 76638
rect 66668 76972 66724 77028
rect 64764 76578 64820 76580
rect 64764 76526 64766 76578
rect 64766 76526 64818 76578
rect 64818 76526 64820 76578
rect 64764 76524 64820 76526
rect 66444 76578 66500 76580
rect 66444 76526 66446 76578
rect 66446 76526 66498 76578
rect 66498 76526 66500 76578
rect 66444 76524 66500 76526
rect 66668 76524 66724 76580
rect 64316 74898 64372 74900
rect 64316 74846 64318 74898
rect 64318 74846 64370 74898
rect 64370 74846 64372 74898
rect 64316 74844 64372 74846
rect 64428 76300 64484 76356
rect 64540 75794 64596 75796
rect 64540 75742 64542 75794
rect 64542 75742 64594 75794
rect 64594 75742 64596 75794
rect 64540 75740 64596 75742
rect 64428 75068 64484 75124
rect 65436 75122 65492 75124
rect 65436 75070 65438 75122
rect 65438 75070 65490 75122
rect 65490 75070 65492 75122
rect 65436 75068 65492 75070
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 66444 75740 66500 75796
rect 67228 76578 67284 76580
rect 67228 76526 67230 76578
rect 67230 76526 67282 76578
rect 67282 76526 67284 76578
rect 67228 76524 67284 76526
rect 66780 76412 66836 76468
rect 66220 75628 66276 75684
rect 66892 76188 66948 76244
rect 67228 75964 67284 76020
rect 66892 75628 66948 75684
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 64428 74172 64484 74228
rect 64092 73500 64148 73556
rect 65324 73554 65380 73556
rect 65324 73502 65326 73554
rect 65326 73502 65378 73554
rect 65378 73502 65380 73554
rect 65324 73500 65380 73502
rect 65548 73500 65604 73556
rect 64764 72940 64820 72996
rect 63980 72156 64036 72212
rect 64428 72268 64484 72324
rect 64204 72156 64260 72212
rect 65324 72156 65380 72212
rect 63196 71650 63252 71652
rect 63196 71598 63198 71650
rect 63198 71598 63250 71650
rect 63250 71598 63252 71650
rect 63196 71596 63252 71598
rect 63756 71596 63812 71652
rect 62860 71036 62916 71092
rect 63308 71036 63364 71092
rect 62972 70364 63028 70420
rect 62412 68348 62468 68404
rect 62524 68012 62580 68068
rect 61628 66274 61684 66276
rect 61628 66222 61630 66274
rect 61630 66222 61682 66274
rect 61682 66222 61684 66274
rect 61628 66220 61684 66222
rect 63196 68626 63252 68628
rect 63196 68574 63198 68626
rect 63198 68574 63250 68626
rect 63250 68574 63252 68626
rect 63196 68572 63252 68574
rect 63196 68348 63252 68404
rect 63644 68796 63700 68852
rect 63420 68012 63476 68068
rect 63532 68572 63588 68628
rect 61852 65548 61908 65604
rect 60508 64764 60564 64820
rect 59836 64706 59892 64708
rect 59836 64654 59838 64706
rect 59838 64654 59890 64706
rect 59890 64654 59892 64706
rect 59836 64652 59892 64654
rect 61740 64818 61796 64820
rect 61740 64766 61742 64818
rect 61742 64766 61794 64818
rect 61794 64766 61796 64818
rect 61740 64764 61796 64766
rect 60284 64482 60340 64484
rect 60284 64430 60286 64482
rect 60286 64430 60338 64482
rect 60338 64430 60340 64482
rect 60284 64428 60340 64430
rect 61740 64428 61796 64484
rect 61628 64316 61684 64372
rect 62860 65548 62916 65604
rect 61964 64204 62020 64260
rect 60396 63756 60452 63812
rect 59276 62748 59332 62804
rect 60060 62524 60116 62580
rect 60284 62748 60340 62804
rect 59164 61458 59220 61460
rect 59164 61406 59166 61458
rect 59166 61406 59218 61458
rect 59218 61406 59220 61458
rect 59164 61404 59220 61406
rect 60172 61458 60228 61460
rect 60172 61406 60174 61458
rect 60174 61406 60226 61458
rect 60226 61406 60228 61458
rect 60172 61404 60228 61406
rect 59276 61292 59332 61348
rect 59724 61346 59780 61348
rect 59724 61294 59726 61346
rect 59726 61294 59778 61346
rect 59778 61294 59780 61346
rect 59724 61292 59780 61294
rect 59724 61068 59780 61124
rect 57372 60732 57428 60788
rect 57260 60226 57316 60228
rect 57260 60174 57262 60226
rect 57262 60174 57314 60226
rect 57314 60174 57316 60226
rect 57260 60172 57316 60174
rect 57260 59890 57316 59892
rect 57260 59838 57262 59890
rect 57262 59838 57314 59890
rect 57314 59838 57316 59890
rect 57260 59836 57316 59838
rect 57372 59724 57428 59780
rect 58044 59836 58100 59892
rect 57596 59330 57652 59332
rect 57596 59278 57598 59330
rect 57598 59278 57650 59330
rect 57650 59278 57652 59330
rect 57596 59276 57652 59278
rect 57708 59218 57764 59220
rect 57708 59166 57710 59218
rect 57710 59166 57762 59218
rect 57762 59166 57764 59218
rect 57708 59164 57764 59166
rect 57260 58828 57316 58884
rect 57596 58604 57652 58660
rect 57932 58940 57988 58996
rect 58380 59890 58436 59892
rect 58380 59838 58382 59890
rect 58382 59838 58434 59890
rect 58434 59838 58436 59890
rect 58380 59836 58436 59838
rect 58492 59724 58548 59780
rect 58156 59612 58212 59668
rect 58492 59500 58548 59556
rect 58156 59442 58212 59444
rect 58156 59390 58158 59442
rect 58158 59390 58210 59442
rect 58210 59390 58212 59442
rect 58156 59388 58212 59390
rect 57260 57708 57316 57764
rect 57372 57820 57428 57876
rect 57372 57596 57428 57652
rect 57708 57762 57764 57764
rect 57708 57710 57710 57762
rect 57710 57710 57762 57762
rect 57762 57710 57764 57762
rect 57708 57708 57764 57710
rect 57484 57036 57540 57092
rect 57484 56866 57540 56868
rect 57484 56814 57486 56866
rect 57486 56814 57538 56866
rect 57538 56814 57540 56866
rect 57484 56812 57540 56814
rect 57372 56754 57428 56756
rect 57372 56702 57374 56754
rect 57374 56702 57426 56754
rect 57426 56702 57428 56754
rect 57372 56700 57428 56702
rect 57596 56364 57652 56420
rect 57372 56306 57428 56308
rect 57372 56254 57374 56306
rect 57374 56254 57426 56306
rect 57426 56254 57428 56306
rect 57372 56252 57428 56254
rect 57036 55244 57092 55300
rect 55692 54460 55748 54516
rect 56028 54236 56084 54292
rect 55356 51660 55412 51716
rect 53900 48466 53956 48468
rect 53900 48414 53902 48466
rect 53902 48414 53954 48466
rect 53954 48414 53956 48466
rect 53900 48412 53956 48414
rect 54124 48354 54180 48356
rect 54124 48302 54126 48354
rect 54126 48302 54178 48354
rect 54178 48302 54180 48354
rect 54124 48300 54180 48302
rect 53676 48188 53732 48244
rect 53564 48076 53620 48132
rect 53340 47068 53396 47124
rect 53676 47068 53732 47124
rect 53676 46844 53732 46900
rect 54236 46898 54292 46900
rect 54236 46846 54238 46898
rect 54238 46846 54290 46898
rect 54290 46846 54292 46898
rect 54236 46844 54292 46846
rect 52332 44098 52388 44100
rect 52332 44046 52334 44098
rect 52334 44046 52386 44098
rect 52386 44046 52388 44098
rect 52332 44044 52388 44046
rect 53228 44044 53284 44100
rect 52780 43650 52836 43652
rect 52780 43598 52782 43650
rect 52782 43598 52834 43650
rect 52834 43598 52836 43650
rect 52780 43596 52836 43598
rect 52220 43484 52276 43540
rect 52332 43260 52388 43316
rect 52668 42028 52724 42084
rect 52444 41858 52500 41860
rect 52444 41806 52446 41858
rect 52446 41806 52498 41858
rect 52498 41806 52500 41858
rect 52444 41804 52500 41806
rect 52556 41244 52612 41300
rect 53452 43484 53508 43540
rect 53340 43260 53396 43316
rect 53452 41858 53508 41860
rect 53452 41806 53454 41858
rect 53454 41806 53506 41858
rect 53506 41806 53508 41858
rect 53452 41804 53508 41806
rect 53116 41132 53172 41188
rect 52332 41074 52388 41076
rect 52332 41022 52334 41074
rect 52334 41022 52386 41074
rect 52386 41022 52388 41074
rect 52332 41020 52388 41022
rect 52332 39452 52388 39508
rect 49196 37324 49252 37380
rect 48972 36652 49028 36708
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50316 37378 50372 37380
rect 50316 37326 50318 37378
rect 50318 37326 50370 37378
rect 50370 37326 50372 37378
rect 50316 37324 50372 37326
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 52668 38162 52724 38164
rect 52668 38110 52670 38162
rect 52670 38110 52722 38162
rect 52722 38110 52724 38162
rect 52668 38108 52724 38110
rect 51436 37100 51492 37156
rect 51100 36706 51156 36708
rect 51100 36654 51102 36706
rect 51102 36654 51154 36706
rect 51154 36654 51156 36706
rect 51100 36652 51156 36654
rect 52444 37154 52500 37156
rect 52444 37102 52446 37154
rect 52446 37102 52498 37154
rect 52498 37102 52500 37154
rect 52444 37100 52500 37102
rect 52220 36482 52276 36484
rect 52220 36430 52222 36482
rect 52222 36430 52274 36482
rect 52274 36430 52276 36482
rect 52220 36428 52276 36430
rect 53452 38780 53508 38836
rect 52892 38668 52948 38724
rect 53452 38162 53508 38164
rect 53452 38110 53454 38162
rect 53454 38110 53506 38162
rect 53506 38110 53508 38162
rect 53452 38108 53508 38110
rect 52780 36428 52836 36484
rect 53340 36482 53396 36484
rect 53340 36430 53342 36482
rect 53342 36430 53394 36482
rect 53394 36430 53396 36482
rect 53340 36428 53396 36430
rect 52108 36370 52164 36372
rect 52108 36318 52110 36370
rect 52110 36318 52162 36370
rect 52162 36318 52164 36370
rect 52108 36316 52164 36318
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 55020 50204 55076 50260
rect 54124 45276 54180 45332
rect 53788 43538 53844 43540
rect 53788 43486 53790 43538
rect 53790 43486 53842 43538
rect 53842 43486 53844 43538
rect 53788 43484 53844 43486
rect 54348 43650 54404 43652
rect 54348 43598 54350 43650
rect 54350 43598 54402 43650
rect 54402 43598 54404 43650
rect 54348 43596 54404 43598
rect 54908 48802 54964 48804
rect 54908 48750 54910 48802
rect 54910 48750 54962 48802
rect 54962 48750 54964 48802
rect 54908 48748 54964 48750
rect 54796 48524 54852 48580
rect 55132 49868 55188 49924
rect 55580 49922 55636 49924
rect 55580 49870 55582 49922
rect 55582 49870 55634 49922
rect 55634 49870 55636 49922
rect 55580 49868 55636 49870
rect 54908 48188 54964 48244
rect 55244 48076 55300 48132
rect 56476 54236 56532 54292
rect 56364 53730 56420 53732
rect 56364 53678 56366 53730
rect 56366 53678 56418 53730
rect 56418 53678 56420 53730
rect 56364 53676 56420 53678
rect 56700 54012 56756 54068
rect 57372 54236 57428 54292
rect 57932 57708 57988 57764
rect 57484 54012 57540 54068
rect 57036 53676 57092 53732
rect 57484 53730 57540 53732
rect 57484 53678 57486 53730
rect 57486 53678 57538 53730
rect 57538 53678 57540 53730
rect 57484 53676 57540 53678
rect 57820 53676 57876 53732
rect 56476 53506 56532 53508
rect 56476 53454 56478 53506
rect 56478 53454 56530 53506
rect 56530 53454 56532 53506
rect 56476 53452 56532 53454
rect 57036 53452 57092 53508
rect 56588 52220 56644 52276
rect 56252 51436 56308 51492
rect 56924 51436 56980 51492
rect 56364 50764 56420 50820
rect 56812 50652 56868 50708
rect 56028 49868 56084 49924
rect 56476 49980 56532 50036
rect 56700 50034 56756 50036
rect 56700 49982 56702 50034
rect 56702 49982 56754 50034
rect 56754 49982 56756 50034
rect 56700 49980 56756 49982
rect 56476 49532 56532 49588
rect 55244 47740 55300 47796
rect 54908 47458 54964 47460
rect 54908 47406 54910 47458
rect 54910 47406 54962 47458
rect 54962 47406 54964 47458
rect 54908 47404 54964 47406
rect 55244 46898 55300 46900
rect 55244 46846 55246 46898
rect 55246 46846 55298 46898
rect 55298 46846 55300 46898
rect 55244 46844 55300 46846
rect 55468 45276 55524 45332
rect 55692 48076 55748 48132
rect 56588 48412 56644 48468
rect 56476 48354 56532 48356
rect 56476 48302 56478 48354
rect 56478 48302 56530 48354
rect 56530 48302 56532 48354
rect 56476 48300 56532 48302
rect 56588 48242 56644 48244
rect 56588 48190 56590 48242
rect 56590 48190 56642 48242
rect 56642 48190 56644 48242
rect 56588 48188 56644 48190
rect 56700 45276 56756 45332
rect 54124 42082 54180 42084
rect 54124 42030 54126 42082
rect 54126 42030 54178 42082
rect 54178 42030 54180 42082
rect 54124 42028 54180 42030
rect 54684 42028 54740 42084
rect 54236 41298 54292 41300
rect 54236 41246 54238 41298
rect 54238 41246 54290 41298
rect 54290 41246 54292 41298
rect 54236 41244 54292 41246
rect 55132 41298 55188 41300
rect 55132 41246 55134 41298
rect 55134 41246 55186 41298
rect 55186 41246 55188 41298
rect 55132 41244 55188 41246
rect 54684 41074 54740 41076
rect 54684 41022 54686 41074
rect 54686 41022 54738 41074
rect 54738 41022 54740 41074
rect 54684 41020 54740 41022
rect 55580 40402 55636 40404
rect 55580 40350 55582 40402
rect 55582 40350 55634 40402
rect 55634 40350 55636 40402
rect 55580 40348 55636 40350
rect 53676 39452 53732 39508
rect 54572 38946 54628 38948
rect 54572 38894 54574 38946
rect 54574 38894 54626 38946
rect 54626 38894 54628 38946
rect 54572 38892 54628 38894
rect 55468 38892 55524 38948
rect 53788 38834 53844 38836
rect 53788 38782 53790 38834
rect 53790 38782 53842 38834
rect 53842 38782 53844 38834
rect 53788 38780 53844 38782
rect 56588 43596 56644 43652
rect 56700 44380 56756 44436
rect 57596 52162 57652 52164
rect 57596 52110 57598 52162
rect 57598 52110 57650 52162
rect 57650 52110 57652 52162
rect 57596 52108 57652 52110
rect 58492 58434 58548 58436
rect 58492 58382 58494 58434
rect 58494 58382 58546 58434
rect 58546 58382 58548 58434
rect 58492 58380 58548 58382
rect 58380 57820 58436 57876
rect 58268 56754 58324 56756
rect 58268 56702 58270 56754
rect 58270 56702 58322 56754
rect 58322 56702 58324 56754
rect 58268 56700 58324 56702
rect 58156 56642 58212 56644
rect 58156 56590 58158 56642
rect 58158 56590 58210 56642
rect 58210 56590 58212 56642
rect 58156 56588 58212 56590
rect 58156 56028 58212 56084
rect 58156 55468 58212 55524
rect 58940 59612 58996 59668
rect 58940 59164 58996 59220
rect 58716 56700 58772 56756
rect 59612 58380 59668 58436
rect 59164 56028 59220 56084
rect 60396 61068 60452 61124
rect 59836 58434 59892 58436
rect 59836 58382 59838 58434
rect 59838 58382 59890 58434
rect 59890 58382 59892 58434
rect 59836 58380 59892 58382
rect 58156 55356 58212 55412
rect 58268 51938 58324 51940
rect 58268 51886 58270 51938
rect 58270 51886 58322 51938
rect 58322 51886 58324 51938
rect 58268 51884 58324 51886
rect 57372 51100 57428 51156
rect 58380 50706 58436 50708
rect 58380 50654 58382 50706
rect 58382 50654 58434 50706
rect 58434 50654 58436 50706
rect 58380 50652 58436 50654
rect 57484 50594 57540 50596
rect 57484 50542 57486 50594
rect 57486 50542 57538 50594
rect 57538 50542 57540 50594
rect 57484 50540 57540 50542
rect 58044 50594 58100 50596
rect 58044 50542 58046 50594
rect 58046 50542 58098 50594
rect 58098 50542 58100 50594
rect 58044 50540 58100 50542
rect 57596 50428 57652 50484
rect 57036 49980 57092 50036
rect 57484 49810 57540 49812
rect 57484 49758 57486 49810
rect 57486 49758 57538 49810
rect 57538 49758 57540 49810
rect 57484 49756 57540 49758
rect 57036 48748 57092 48804
rect 57484 49532 57540 49588
rect 57372 48354 57428 48356
rect 57372 48302 57374 48354
rect 57374 48302 57426 48354
rect 57426 48302 57428 48354
rect 57372 48300 57428 48302
rect 57596 48748 57652 48804
rect 58156 49532 58212 49588
rect 58380 48188 58436 48244
rect 57708 48076 57764 48132
rect 59276 54236 59332 54292
rect 58716 51548 58772 51604
rect 58940 51884 58996 51940
rect 58716 51324 58772 51380
rect 58716 50428 58772 50484
rect 58604 49756 58660 49812
rect 58604 49196 58660 49252
rect 58828 50764 58884 50820
rect 58604 48466 58660 48468
rect 58604 48414 58606 48466
rect 58606 48414 58658 48466
rect 58658 48414 58660 48466
rect 58604 48412 58660 48414
rect 58268 47068 58324 47124
rect 58156 44492 58212 44548
rect 56476 41970 56532 41972
rect 56476 41918 56478 41970
rect 56478 41918 56530 41970
rect 56530 41918 56532 41970
rect 56476 41916 56532 41918
rect 56028 40402 56084 40404
rect 56028 40350 56030 40402
rect 56030 40350 56082 40402
rect 56082 40350 56084 40402
rect 56028 40348 56084 40350
rect 57036 41916 57092 41972
rect 56924 41804 56980 41860
rect 56924 41356 56980 41412
rect 57036 40348 57092 40404
rect 54348 36540 54404 36596
rect 53676 36316 53732 36372
rect 54124 36428 54180 36484
rect 55580 36540 55636 36596
rect 55692 37826 55748 37828
rect 55692 37774 55694 37826
rect 55694 37774 55746 37826
rect 55746 37774 55748 37826
rect 55692 37772 55748 37774
rect 54124 35868 54180 35924
rect 52892 35644 52948 35700
rect 49868 34914 49924 34916
rect 49868 34862 49870 34914
rect 49870 34862 49922 34914
rect 49922 34862 49924 34914
rect 49868 34860 49924 34862
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 53564 35644 53620 35700
rect 51324 35420 51380 35476
rect 52668 35308 52724 35364
rect 53564 35474 53620 35476
rect 53564 35422 53566 35474
rect 53566 35422 53618 35474
rect 53618 35422 53620 35474
rect 53564 35420 53620 35422
rect 53900 35308 53956 35364
rect 53676 34860 53732 34916
rect 53004 34748 53060 34804
rect 54012 34748 54068 34804
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 53116 33404 53172 33460
rect 53900 34130 53956 34132
rect 53900 34078 53902 34130
rect 53902 34078 53954 34130
rect 53954 34078 53956 34130
rect 53900 34076 53956 34078
rect 53788 33458 53844 33460
rect 53788 33406 53790 33458
rect 53790 33406 53842 33458
rect 53842 33406 53844 33458
rect 53788 33404 53844 33406
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 55244 35922 55300 35924
rect 55244 35870 55246 35922
rect 55246 35870 55298 35922
rect 55298 35870 55300 35922
rect 55244 35868 55300 35870
rect 54460 35644 54516 35700
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 14252 3276 14308 3332
rect 19404 3330 19460 3332
rect 19404 3278 19406 3330
rect 19406 3278 19458 3330
rect 19458 3278 19460 3330
rect 19404 3276 19460 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 43708 3388 43764 3444
rect 31836 2828 31892 2884
rect 44268 3442 44324 3444
rect 44268 3390 44270 3442
rect 44270 3390 44322 3442
rect 44322 3390 44324 3442
rect 44268 3388 44324 3390
rect 44940 3442 44996 3444
rect 44940 3390 44942 3442
rect 44942 3390 44994 3442
rect 44994 3390 44996 3442
rect 44940 3388 44996 3390
rect 54684 34802 54740 34804
rect 54684 34750 54686 34802
rect 54686 34750 54738 34802
rect 54738 34750 54740 34802
rect 54684 34748 54740 34750
rect 56476 37266 56532 37268
rect 56476 37214 56478 37266
rect 56478 37214 56530 37266
rect 56530 37214 56532 37266
rect 56476 37212 56532 37214
rect 55692 34748 55748 34804
rect 57260 37772 57316 37828
rect 57372 37660 57428 37716
rect 56700 34972 56756 35028
rect 57596 43650 57652 43652
rect 57596 43598 57598 43650
rect 57598 43598 57650 43650
rect 57650 43598 57652 43650
rect 57596 43596 57652 43598
rect 57932 42812 57988 42868
rect 57596 41916 57652 41972
rect 57708 41186 57764 41188
rect 57708 41134 57710 41186
rect 57710 41134 57762 41186
rect 57762 41134 57764 41186
rect 57708 41132 57764 41134
rect 58156 40908 58212 40964
rect 58156 37772 58212 37828
rect 58044 37660 58100 37716
rect 57708 37266 57764 37268
rect 57708 37214 57710 37266
rect 57710 37214 57762 37266
rect 57762 37214 57764 37266
rect 57708 37212 57764 37214
rect 57484 35420 57540 35476
rect 57372 35026 57428 35028
rect 57372 34974 57374 35026
rect 57374 34974 57426 35026
rect 57426 34974 57428 35026
rect 57372 34972 57428 34974
rect 56700 34188 56756 34244
rect 54460 34076 54516 34132
rect 56700 34018 56756 34020
rect 56700 33966 56702 34018
rect 56702 33966 56754 34018
rect 56754 33966 56756 34018
rect 56700 33964 56756 33966
rect 54796 32562 54852 32564
rect 54796 32510 54798 32562
rect 54798 32510 54850 32562
rect 54850 32510 54852 32562
rect 54796 32508 54852 32510
rect 56476 33180 56532 33236
rect 55916 33068 55972 33124
rect 55468 32562 55524 32564
rect 55468 32510 55470 32562
rect 55470 32510 55522 32562
rect 55522 32510 55524 32562
rect 55468 32508 55524 32510
rect 55804 32562 55860 32564
rect 55804 32510 55806 32562
rect 55806 32510 55858 32562
rect 55858 32510 55860 32562
rect 55804 32508 55860 32510
rect 57372 33292 57428 33348
rect 57036 33180 57092 33236
rect 57372 32508 57428 32564
rect 58044 35810 58100 35812
rect 58044 35758 58046 35810
rect 58046 35758 58098 35810
rect 58098 35758 58100 35810
rect 58044 35756 58100 35758
rect 58156 35420 58212 35476
rect 58268 34076 58324 34132
rect 57932 33964 57988 34020
rect 57820 32786 57876 32788
rect 57820 32734 57822 32786
rect 57822 32734 57874 32786
rect 57874 32734 57876 32786
rect 57820 32732 57876 32734
rect 58044 33122 58100 33124
rect 58044 33070 58046 33122
rect 58046 33070 58098 33122
rect 58098 33070 58100 33122
rect 58044 33068 58100 33070
rect 58492 44492 58548 44548
rect 59388 51436 59444 51492
rect 59164 50988 59220 51044
rect 58940 50540 58996 50596
rect 58940 48242 58996 48244
rect 58940 48190 58942 48242
rect 58942 48190 58994 48242
rect 58994 48190 58996 48242
rect 58940 48188 58996 48190
rect 59276 47740 59332 47796
rect 59052 47068 59108 47124
rect 59500 47068 59556 47124
rect 58828 44492 58884 44548
rect 59276 44492 59332 44548
rect 58604 44434 58660 44436
rect 58604 44382 58606 44434
rect 58606 44382 58658 44434
rect 58658 44382 58660 44434
rect 58604 44380 58660 44382
rect 59724 54738 59780 54740
rect 59724 54686 59726 54738
rect 59726 54686 59778 54738
rect 59778 54686 59780 54738
rect 59724 54684 59780 54686
rect 59948 54236 60004 54292
rect 60396 60620 60452 60676
rect 61180 63922 61236 63924
rect 61180 63870 61182 63922
rect 61182 63870 61234 63922
rect 61234 63870 61236 63922
rect 61180 63868 61236 63870
rect 61852 61852 61908 61908
rect 62188 62914 62244 62916
rect 62188 62862 62190 62914
rect 62190 62862 62242 62914
rect 62242 62862 62244 62914
rect 62188 62860 62244 62862
rect 62188 62466 62244 62468
rect 62188 62414 62190 62466
rect 62190 62414 62242 62466
rect 62242 62414 62244 62466
rect 62188 62412 62244 62414
rect 63308 62578 63364 62580
rect 63308 62526 63310 62578
rect 63310 62526 63362 62578
rect 63362 62526 63364 62578
rect 63308 62524 63364 62526
rect 63196 62466 63252 62468
rect 63196 62414 63198 62466
rect 63198 62414 63250 62466
rect 63250 62414 63252 62466
rect 63196 62412 63252 62414
rect 61628 61292 61684 61348
rect 60508 59836 60564 59892
rect 61068 59388 61124 59444
rect 60956 58380 61012 58436
rect 60620 58322 60676 58324
rect 60620 58270 60622 58322
rect 60622 58270 60674 58322
rect 60674 58270 60676 58322
rect 60620 58268 60676 58270
rect 60396 57036 60452 57092
rect 60284 52892 60340 52948
rect 59724 51490 59780 51492
rect 59724 51438 59726 51490
rect 59726 51438 59778 51490
rect 59778 51438 59780 51490
rect 59724 51436 59780 51438
rect 60284 51378 60340 51380
rect 60284 51326 60286 51378
rect 60286 51326 60338 51378
rect 60338 51326 60340 51378
rect 60284 51324 60340 51326
rect 59724 50764 59780 50820
rect 60172 50706 60228 50708
rect 60172 50654 60174 50706
rect 60174 50654 60226 50706
rect 60226 50654 60228 50706
rect 60172 50652 60228 50654
rect 59724 48130 59780 48132
rect 59724 48078 59726 48130
rect 59726 48078 59778 48130
rect 59778 48078 59780 48130
rect 59724 48076 59780 48078
rect 59948 47570 60004 47572
rect 59948 47518 59950 47570
rect 59950 47518 60002 47570
rect 60002 47518 60004 47570
rect 59948 47516 60004 47518
rect 59612 43820 59668 43876
rect 58716 43372 58772 43428
rect 59276 43426 59332 43428
rect 59276 43374 59278 43426
rect 59278 43374 59330 43426
rect 59330 43374 59332 43426
rect 59276 43372 59332 43374
rect 58940 42812 58996 42868
rect 58604 41186 58660 41188
rect 58604 41134 58606 41186
rect 58606 41134 58658 41186
rect 58658 41134 58660 41186
rect 58604 41132 58660 41134
rect 59500 40908 59556 40964
rect 60620 57036 60676 57092
rect 60620 55468 60676 55524
rect 60508 55020 60564 55076
rect 61852 60844 61908 60900
rect 62860 61852 62916 61908
rect 62748 61628 62804 61684
rect 63420 62412 63476 62468
rect 62972 61516 63028 61572
rect 62300 60844 62356 60900
rect 61740 59388 61796 59444
rect 61404 57820 61460 57876
rect 60844 55132 60900 55188
rect 61180 55356 61236 55412
rect 60956 53788 61012 53844
rect 61068 54460 61124 54516
rect 60844 53116 60900 53172
rect 61292 55186 61348 55188
rect 61292 55134 61294 55186
rect 61294 55134 61346 55186
rect 61346 55134 61348 55186
rect 61292 55132 61348 55134
rect 61516 55132 61572 55188
rect 61404 54626 61460 54628
rect 61404 54574 61406 54626
rect 61406 54574 61458 54626
rect 61458 54574 61460 54626
rect 61404 54572 61460 54574
rect 60844 51884 60900 51940
rect 60844 51378 60900 51380
rect 60844 51326 60846 51378
rect 60846 51326 60898 51378
rect 60898 51326 60900 51378
rect 60844 51324 60900 51326
rect 61180 51266 61236 51268
rect 61180 51214 61182 51266
rect 61182 51214 61234 51266
rect 61234 51214 61236 51266
rect 61180 51212 61236 51214
rect 60620 48802 60676 48804
rect 60620 48750 60622 48802
rect 60622 48750 60674 48802
rect 60674 48750 60676 48802
rect 60620 48748 60676 48750
rect 60620 48242 60676 48244
rect 60620 48190 60622 48242
rect 60622 48190 60674 48242
rect 60674 48190 60676 48242
rect 60620 48188 60676 48190
rect 60844 47964 60900 48020
rect 60620 47404 60676 47460
rect 60956 46732 61012 46788
rect 61068 47292 61124 47348
rect 60396 43260 60452 43316
rect 60396 42866 60452 42868
rect 60396 42814 60398 42866
rect 60398 42814 60450 42866
rect 60450 42814 60452 42866
rect 60396 42812 60452 42814
rect 60172 41804 60228 41860
rect 60732 41916 60788 41972
rect 58940 40402 58996 40404
rect 58940 40350 58942 40402
rect 58942 40350 58994 40402
rect 58994 40350 58996 40402
rect 58940 40348 58996 40350
rect 60732 39564 60788 39620
rect 60284 39340 60340 39396
rect 59948 39004 60004 39060
rect 61068 38108 61124 38164
rect 58716 37660 58772 37716
rect 59388 37660 59444 37716
rect 58828 37436 58884 37492
rect 59724 37660 59780 37716
rect 59836 37490 59892 37492
rect 59836 37438 59838 37490
rect 59838 37438 59890 37490
rect 59890 37438 59892 37490
rect 59836 37436 59892 37438
rect 58604 35756 58660 35812
rect 58380 33964 58436 34020
rect 58716 35474 58772 35476
rect 58716 35422 58718 35474
rect 58718 35422 58770 35474
rect 58770 35422 58772 35474
rect 58716 35420 58772 35422
rect 60284 35698 60340 35700
rect 60284 35646 60286 35698
rect 60286 35646 60338 35698
rect 60338 35646 60340 35698
rect 60284 35644 60340 35646
rect 59948 34636 60004 34692
rect 58380 33346 58436 33348
rect 58380 33294 58382 33346
rect 58382 33294 58434 33346
rect 58434 33294 58436 33346
rect 58380 33292 58436 33294
rect 61628 52220 61684 52276
rect 61628 51324 61684 51380
rect 65324 71596 65380 71652
rect 65436 72268 65492 72324
rect 64316 71090 64372 71092
rect 64316 71038 64318 71090
rect 64318 71038 64370 71090
rect 64370 71038 64372 71090
rect 64316 71036 64372 71038
rect 63868 70418 63924 70420
rect 63868 70366 63870 70418
rect 63870 70366 63922 70418
rect 63922 70366 63924 70418
rect 63868 70364 63924 70366
rect 64764 70364 64820 70420
rect 63868 68626 63924 68628
rect 63868 68574 63870 68626
rect 63870 68574 63922 68626
rect 63922 68574 63924 68626
rect 63868 68572 63924 68574
rect 63756 68012 63812 68068
rect 64316 68012 64372 68068
rect 64988 65660 65044 65716
rect 64316 65602 64372 65604
rect 64316 65550 64318 65602
rect 64318 65550 64370 65602
rect 64370 65550 64372 65602
rect 64316 65548 64372 65550
rect 64092 64706 64148 64708
rect 64092 64654 64094 64706
rect 64094 64654 64146 64706
rect 64146 64654 64148 64706
rect 64092 64652 64148 64654
rect 63980 62578 64036 62580
rect 63980 62526 63982 62578
rect 63982 62526 64034 62578
rect 64034 62526 64036 62578
rect 63980 62524 64036 62526
rect 64876 62188 64932 62244
rect 63756 61628 63812 61684
rect 63644 61068 63700 61124
rect 63532 60508 63588 60564
rect 63644 60060 63700 60116
rect 63084 59948 63140 60004
rect 61852 59052 61908 59108
rect 62412 59106 62468 59108
rect 62412 59054 62414 59106
rect 62414 59054 62466 59106
rect 62466 59054 62468 59106
rect 62412 59052 62468 59054
rect 62748 58940 62804 58996
rect 62412 55356 62468 55412
rect 62412 55020 62468 55076
rect 62300 54684 62356 54740
rect 62076 54572 62132 54628
rect 61852 54460 61908 54516
rect 62188 53788 62244 53844
rect 61964 52946 62020 52948
rect 61964 52894 61966 52946
rect 61966 52894 62018 52946
rect 62018 52894 62020 52946
rect 61964 52892 62020 52894
rect 62524 52946 62580 52948
rect 62524 52894 62526 52946
rect 62526 52894 62578 52946
rect 62578 52894 62580 52946
rect 62524 52892 62580 52894
rect 62076 52332 62132 52388
rect 62076 51436 62132 51492
rect 61740 51100 61796 51156
rect 61404 47516 61460 47572
rect 61852 48860 61908 48916
rect 61516 47404 61572 47460
rect 61404 47346 61460 47348
rect 61404 47294 61406 47346
rect 61406 47294 61458 47346
rect 61458 47294 61460 47346
rect 61404 47292 61460 47294
rect 61964 49868 62020 49924
rect 61740 48412 61796 48468
rect 62636 52162 62692 52164
rect 62636 52110 62638 52162
rect 62638 52110 62690 52162
rect 62690 52110 62692 52162
rect 62636 52108 62692 52110
rect 62188 48748 62244 48804
rect 62412 50988 62468 51044
rect 61852 48018 61908 48020
rect 61852 47966 61854 48018
rect 61854 47966 61906 48018
rect 61906 47966 61908 48018
rect 61852 47964 61908 47966
rect 61852 47516 61908 47572
rect 61404 44994 61460 44996
rect 61404 44942 61406 44994
rect 61406 44942 61458 44994
rect 61458 44942 61460 44994
rect 61404 44940 61460 44942
rect 62300 47964 62356 48020
rect 61964 47292 62020 47348
rect 62188 46786 62244 46788
rect 62188 46734 62190 46786
rect 62190 46734 62242 46786
rect 62242 46734 62244 46786
rect 62188 46732 62244 46734
rect 61852 44156 61908 44212
rect 61292 41916 61348 41972
rect 61852 41916 61908 41972
rect 62076 43260 62132 43316
rect 62636 50482 62692 50484
rect 62636 50430 62638 50482
rect 62638 50430 62690 50482
rect 62690 50430 62692 50482
rect 62636 50428 62692 50430
rect 62524 49810 62580 49812
rect 62524 49758 62526 49810
rect 62526 49758 62578 49810
rect 62578 49758 62580 49810
rect 62524 49756 62580 49758
rect 62636 48748 62692 48804
rect 62524 48524 62580 48580
rect 63196 58604 63252 58660
rect 63084 54684 63140 54740
rect 62860 54572 62916 54628
rect 63196 53170 63252 53172
rect 63196 53118 63198 53170
rect 63198 53118 63250 53170
rect 63250 53118 63252 53170
rect 63196 53116 63252 53118
rect 62972 51266 63028 51268
rect 62972 51214 62974 51266
rect 62974 51214 63026 51266
rect 63026 51214 63028 51266
rect 62972 51212 63028 51214
rect 62748 48636 62804 48692
rect 63196 50428 63252 50484
rect 62860 48354 62916 48356
rect 62860 48302 62862 48354
rect 62862 48302 62914 48354
rect 62914 48302 62916 48354
rect 62860 48300 62916 48302
rect 62524 47292 62580 47348
rect 62524 43708 62580 43764
rect 61740 41692 61796 41748
rect 61292 40348 61348 40404
rect 62748 42812 62804 42868
rect 62412 41692 62468 41748
rect 62188 41298 62244 41300
rect 62188 41246 62190 41298
rect 62190 41246 62242 41298
rect 62242 41246 62244 41298
rect 62188 41244 62244 41246
rect 63084 41132 63140 41188
rect 62748 41020 62804 41076
rect 62188 40626 62244 40628
rect 62188 40574 62190 40626
rect 62190 40574 62242 40626
rect 62242 40574 62244 40626
rect 62188 40572 62244 40574
rect 63084 40572 63140 40628
rect 62748 40460 62804 40516
rect 61740 39618 61796 39620
rect 61740 39566 61742 39618
rect 61742 39566 61794 39618
rect 61794 39566 61796 39618
rect 61740 39564 61796 39566
rect 61516 38722 61572 38724
rect 61516 38670 61518 38722
rect 61518 38670 61570 38722
rect 61570 38670 61572 38722
rect 61516 38668 61572 38670
rect 61516 38162 61572 38164
rect 61516 38110 61518 38162
rect 61518 38110 61570 38162
rect 61570 38110 61572 38162
rect 61516 38108 61572 38110
rect 61292 37996 61348 38052
rect 61180 37436 61236 37492
rect 61068 35756 61124 35812
rect 60620 34972 60676 35028
rect 61516 37772 61572 37828
rect 61516 36988 61572 37044
rect 62300 39618 62356 39620
rect 62300 39566 62302 39618
rect 62302 39566 62354 39618
rect 62354 39566 62356 39618
rect 62300 39564 62356 39566
rect 62524 39340 62580 39396
rect 62188 39058 62244 39060
rect 62188 39006 62190 39058
rect 62190 39006 62242 39058
rect 62242 39006 62244 39058
rect 62188 39004 62244 39006
rect 63196 39228 63252 39284
rect 62524 38668 62580 38724
rect 62860 38892 62916 38948
rect 63196 38668 63252 38724
rect 63084 38108 63140 38164
rect 62188 38050 62244 38052
rect 62188 37998 62190 38050
rect 62190 37998 62242 38050
rect 62242 37998 62244 38050
rect 62188 37996 62244 37998
rect 61964 36988 62020 37044
rect 62748 35980 62804 36036
rect 61740 35532 61796 35588
rect 60284 34130 60340 34132
rect 60284 34078 60286 34130
rect 60286 34078 60338 34130
rect 60338 34078 60340 34130
rect 60284 34076 60340 34078
rect 60732 34076 60788 34132
rect 59164 33346 59220 33348
rect 59164 33294 59166 33346
rect 59166 33294 59218 33346
rect 59218 33294 59220 33346
rect 59164 33292 59220 33294
rect 59724 33292 59780 33348
rect 58940 32732 58996 32788
rect 59724 32786 59780 32788
rect 59724 32734 59726 32786
rect 59726 32734 59778 32786
rect 59778 32734 59780 32786
rect 59724 32732 59780 32734
rect 60620 33234 60676 33236
rect 60620 33182 60622 33234
rect 60622 33182 60674 33234
rect 60674 33182 60676 33234
rect 60620 33180 60676 33182
rect 60396 32732 60452 32788
rect 60956 34130 61012 34132
rect 60956 34078 60958 34130
rect 60958 34078 61010 34130
rect 61010 34078 61012 34130
rect 60956 34076 61012 34078
rect 62188 35026 62244 35028
rect 62188 34974 62190 35026
rect 62190 34974 62242 35026
rect 62242 34974 62244 35026
rect 62188 34972 62244 34974
rect 63084 35698 63140 35700
rect 63084 35646 63086 35698
rect 63086 35646 63138 35698
rect 63138 35646 63140 35698
rect 63084 35644 63140 35646
rect 62524 34972 62580 35028
rect 62188 34300 62244 34356
rect 61740 33180 61796 33236
rect 61964 33964 62020 34020
rect 61740 32786 61796 32788
rect 61740 32734 61742 32786
rect 61742 32734 61794 32786
rect 61794 32734 61796 32786
rect 61740 32732 61796 32734
rect 61404 32620 61460 32676
rect 63532 58940 63588 58996
rect 63532 56140 63588 56196
rect 63420 53170 63476 53172
rect 63420 53118 63422 53170
rect 63422 53118 63474 53170
rect 63474 53118 63476 53170
rect 63420 53116 63476 53118
rect 63532 53058 63588 53060
rect 63532 53006 63534 53058
rect 63534 53006 63586 53058
rect 63586 53006 63588 53058
rect 63532 53004 63588 53006
rect 63980 60620 64036 60676
rect 64092 60956 64148 61012
rect 63868 59442 63924 59444
rect 63868 59390 63870 59442
rect 63870 59390 63922 59442
rect 63922 59390 63924 59442
rect 63868 59388 63924 59390
rect 63980 59218 64036 59220
rect 63980 59166 63982 59218
rect 63982 59166 64034 59218
rect 64034 59166 64036 59218
rect 63980 59164 64036 59166
rect 63980 55356 64036 55412
rect 63868 55186 63924 55188
rect 63868 55134 63870 55186
rect 63870 55134 63922 55186
rect 63922 55134 63924 55186
rect 63868 55132 63924 55134
rect 63980 52108 64036 52164
rect 63756 51884 63812 51940
rect 64540 60786 64596 60788
rect 64540 60734 64542 60786
rect 64542 60734 64594 60786
rect 64594 60734 64596 60786
rect 64540 60732 64596 60734
rect 64428 60002 64484 60004
rect 64428 59950 64430 60002
rect 64430 59950 64482 60002
rect 64482 59950 64484 60002
rect 64428 59948 64484 59950
rect 65324 70252 65380 70308
rect 65436 69410 65492 69412
rect 65436 69358 65438 69410
rect 65438 69358 65490 69410
rect 65490 69358 65492 69410
rect 65436 69356 65492 69358
rect 65436 68908 65492 68964
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 65772 72322 65828 72324
rect 65772 72270 65774 72322
rect 65774 72270 65826 72322
rect 65826 72270 65828 72322
rect 65772 72268 65828 72270
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 67340 75852 67396 75908
rect 66332 70700 66388 70756
rect 66780 70306 66836 70308
rect 66780 70254 66782 70306
rect 66782 70254 66834 70306
rect 66834 70254 66836 70306
rect 66780 70252 66836 70254
rect 68572 80220 68628 80276
rect 68236 80108 68292 80164
rect 70476 88844 70532 88900
rect 71596 88898 71652 88900
rect 71596 88846 71598 88898
rect 71598 88846 71650 88898
rect 71650 88846 71652 88898
rect 71596 88844 71652 88846
rect 69804 86658 69860 86660
rect 69804 86606 69806 86658
rect 69806 86606 69858 86658
rect 69858 86606 69860 86658
rect 69804 86604 69860 86606
rect 70252 86604 70308 86660
rect 69468 86434 69524 86436
rect 69468 86382 69470 86434
rect 69470 86382 69522 86434
rect 69522 86382 69524 86434
rect 69468 86380 69524 86382
rect 70364 86380 70420 86436
rect 70140 86268 70196 86324
rect 70364 86044 70420 86100
rect 69468 85762 69524 85764
rect 69468 85710 69470 85762
rect 69470 85710 69522 85762
rect 69522 85710 69524 85762
rect 69468 85708 69524 85710
rect 69244 82236 69300 82292
rect 71932 87836 71988 87892
rect 70588 86380 70644 86436
rect 70700 86268 70756 86324
rect 71932 87388 71988 87444
rect 70476 85708 70532 85764
rect 71372 86546 71428 86548
rect 71372 86494 71374 86546
rect 71374 86494 71426 86546
rect 71426 86494 71428 86546
rect 71372 86492 71428 86494
rect 71036 86380 71092 86436
rect 71596 86044 71652 86100
rect 71708 86658 71764 86660
rect 71708 86606 71710 86658
rect 71710 86606 71762 86658
rect 71762 86606 71764 86658
rect 71708 86604 71764 86606
rect 72492 87276 72548 87332
rect 73164 87388 73220 87444
rect 73724 87330 73780 87332
rect 73724 87278 73726 87330
rect 73726 87278 73778 87330
rect 73778 87278 73780 87330
rect 73724 87276 73780 87278
rect 71260 83244 71316 83300
rect 71596 83298 71652 83300
rect 71596 83246 71598 83298
rect 71598 83246 71650 83298
rect 71650 83246 71652 83298
rect 71596 83244 71652 83246
rect 69468 81340 69524 81396
rect 69244 80556 69300 80612
rect 69468 80274 69524 80276
rect 69468 80222 69470 80274
rect 69470 80222 69522 80274
rect 69522 80222 69524 80274
rect 69468 80220 69524 80222
rect 69692 81394 69748 81396
rect 69692 81342 69694 81394
rect 69694 81342 69746 81394
rect 69746 81342 69748 81394
rect 69692 81340 69748 81342
rect 69244 80162 69300 80164
rect 69244 80110 69246 80162
rect 69246 80110 69298 80162
rect 69298 80110 69300 80162
rect 69244 80108 69300 80110
rect 69580 79996 69636 80052
rect 69580 79772 69636 79828
rect 69692 80892 69748 80948
rect 67676 78316 67732 78372
rect 67788 78706 67844 78708
rect 67788 78654 67790 78706
rect 67790 78654 67842 78706
rect 67842 78654 67844 78706
rect 67788 78652 67844 78654
rect 67788 78204 67844 78260
rect 69020 78652 69076 78708
rect 68124 78204 68180 78260
rect 68460 77420 68516 77476
rect 67900 77250 67956 77252
rect 67900 77198 67902 77250
rect 67902 77198 67954 77250
rect 67954 77198 67956 77250
rect 67900 77196 67956 77198
rect 67788 76636 67844 76692
rect 68124 76466 68180 76468
rect 68124 76414 68126 76466
rect 68126 76414 68178 76466
rect 68178 76414 68180 76466
rect 68124 76412 68180 76414
rect 67788 75964 67844 76020
rect 69356 78540 69412 78596
rect 69804 78764 69860 78820
rect 69580 77196 69636 77252
rect 68012 75682 68068 75684
rect 68012 75630 68014 75682
rect 68014 75630 68066 75682
rect 68066 75630 68068 75682
rect 68012 75628 68068 75630
rect 67564 73500 67620 73556
rect 68124 71036 68180 71092
rect 67452 70476 67508 70532
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 67788 70252 67844 70308
rect 68236 70700 68292 70756
rect 67676 69468 67732 69524
rect 67340 69132 67396 69188
rect 67228 68236 67284 68292
rect 66892 67788 66948 67844
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 65436 65660 65492 65716
rect 65660 65548 65716 65604
rect 66556 66274 66612 66276
rect 66556 66222 66558 66274
rect 66558 66222 66610 66274
rect 66610 66222 66612 66274
rect 66556 66220 66612 66222
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 66332 64652 66388 64708
rect 66220 64146 66276 64148
rect 66220 64094 66222 64146
rect 66222 64094 66274 64146
rect 66274 64094 66276 64146
rect 66220 64092 66276 64094
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 66220 63308 66276 63364
rect 65884 62914 65940 62916
rect 65884 62862 65886 62914
rect 65886 62862 65938 62914
rect 65938 62862 65940 62914
rect 65884 62860 65940 62862
rect 66668 65436 66724 65492
rect 65772 62242 65828 62244
rect 65772 62190 65774 62242
rect 65774 62190 65826 62242
rect 65826 62190 65828 62242
rect 65772 62188 65828 62190
rect 64876 60508 64932 60564
rect 65324 60898 65380 60900
rect 65324 60846 65326 60898
rect 65326 60846 65378 60898
rect 65378 60846 65380 60898
rect 65324 60844 65380 60846
rect 65100 59836 65156 59892
rect 64204 58434 64260 58436
rect 64204 58382 64206 58434
rect 64206 58382 64258 58434
rect 64258 58382 64260 58434
rect 64204 58380 64260 58382
rect 64316 58156 64372 58212
rect 64316 54684 64372 54740
rect 64204 54626 64260 54628
rect 64204 54574 64206 54626
rect 64206 54574 64258 54626
rect 64258 54574 64260 54626
rect 64204 54572 64260 54574
rect 64316 53116 64372 53172
rect 64092 51548 64148 51604
rect 64092 51378 64148 51380
rect 64092 51326 64094 51378
rect 64094 51326 64146 51378
rect 64146 51326 64148 51378
rect 64092 51324 64148 51326
rect 64204 48466 64260 48468
rect 64204 48414 64206 48466
rect 64206 48414 64258 48466
rect 64258 48414 64260 48466
rect 64204 48412 64260 48414
rect 64316 48242 64372 48244
rect 64316 48190 64318 48242
rect 64318 48190 64370 48242
rect 64370 48190 64372 48242
rect 64316 48188 64372 48190
rect 63420 48076 63476 48132
rect 64204 48018 64260 48020
rect 64204 47966 64206 48018
rect 64206 47966 64258 48018
rect 64258 47966 64260 48018
rect 64204 47964 64260 47966
rect 64204 47068 64260 47124
rect 64316 46732 64372 46788
rect 63532 45388 63588 45444
rect 63420 43762 63476 43764
rect 63420 43710 63422 43762
rect 63422 43710 63474 43762
rect 63474 43710 63476 43762
rect 63420 43708 63476 43710
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65996 61682 66052 61684
rect 65996 61630 65998 61682
rect 65998 61630 66050 61682
rect 66050 61630 66052 61682
rect 65996 61628 66052 61630
rect 65548 60844 65604 60900
rect 66220 61068 66276 61124
rect 65884 60732 65940 60788
rect 66668 63868 66724 63924
rect 67004 65772 67060 65828
rect 66556 63308 66612 63364
rect 66556 61628 66612 61684
rect 66668 61010 66724 61012
rect 66668 60958 66670 61010
rect 66670 60958 66722 61010
rect 66722 60958 66724 61010
rect 66668 60956 66724 60958
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65548 59724 65604 59780
rect 65436 59500 65492 59556
rect 65324 59164 65380 59220
rect 64988 58658 65044 58660
rect 64988 58606 64990 58658
rect 64990 58606 65042 58658
rect 65042 58606 65044 58658
rect 64988 58604 65044 58606
rect 64540 58380 64596 58436
rect 64540 53788 64596 53844
rect 65100 58434 65156 58436
rect 65100 58382 65102 58434
rect 65102 58382 65154 58434
rect 65154 58382 65156 58434
rect 65100 58380 65156 58382
rect 64988 58210 65044 58212
rect 64988 58158 64990 58210
rect 64990 58158 65042 58210
rect 65042 58158 65044 58210
rect 64988 58156 65044 58158
rect 65548 58322 65604 58324
rect 65548 58270 65550 58322
rect 65550 58270 65602 58322
rect 65602 58270 65604 58322
rect 65548 58268 65604 58270
rect 66332 59778 66388 59780
rect 66332 59726 66334 59778
rect 66334 59726 66386 59778
rect 66386 59726 66388 59778
rect 66332 59724 66388 59726
rect 67004 63980 67060 64036
rect 66892 62860 66948 62916
rect 67116 62914 67172 62916
rect 67116 62862 67118 62914
rect 67118 62862 67170 62914
rect 67170 62862 67172 62914
rect 67116 62860 67172 62862
rect 67564 68460 67620 68516
rect 67452 67842 67508 67844
rect 67452 67790 67454 67842
rect 67454 67790 67506 67842
rect 67506 67790 67508 67842
rect 67452 67788 67508 67790
rect 68236 69186 68292 69188
rect 68236 69134 68238 69186
rect 68238 69134 68290 69186
rect 68290 69134 68292 69186
rect 68236 69132 68292 69134
rect 68572 73948 68628 74004
rect 69468 74002 69524 74004
rect 69468 73950 69470 74002
rect 69470 73950 69522 74002
rect 69522 73950 69524 74002
rect 69468 73948 69524 73950
rect 70140 81058 70196 81060
rect 70140 81006 70142 81058
rect 70142 81006 70194 81058
rect 70194 81006 70196 81058
rect 70140 81004 70196 81006
rect 71484 81170 71540 81172
rect 71484 81118 71486 81170
rect 71486 81118 71538 81170
rect 71538 81118 71540 81170
rect 71484 81116 71540 81118
rect 70588 80892 70644 80948
rect 70476 80556 70532 80612
rect 70028 80386 70084 80388
rect 70028 80334 70030 80386
rect 70030 80334 70082 80386
rect 70082 80334 70084 80386
rect 70028 80332 70084 80334
rect 70364 80386 70420 80388
rect 70364 80334 70366 80386
rect 70366 80334 70418 80386
rect 70418 80334 70420 80386
rect 70364 80332 70420 80334
rect 70140 80108 70196 80164
rect 70028 78258 70084 78260
rect 70028 78206 70030 78258
rect 70030 78206 70082 78258
rect 70082 78206 70084 78258
rect 70028 78204 70084 78206
rect 70252 79660 70308 79716
rect 70364 80108 70420 80164
rect 70700 80444 70756 80500
rect 71372 80332 71428 80388
rect 70812 80274 70868 80276
rect 70812 80222 70814 80274
rect 70814 80222 70866 80274
rect 70866 80222 70868 80274
rect 70812 80220 70868 80222
rect 70588 78540 70644 78596
rect 71484 80220 71540 80276
rect 71484 79548 71540 79604
rect 71932 86268 71988 86324
rect 73388 86604 73444 86660
rect 72716 86098 72772 86100
rect 72716 86046 72718 86098
rect 72718 86046 72770 86098
rect 72770 86046 72772 86098
rect 72716 86044 72772 86046
rect 73724 86658 73780 86660
rect 73724 86606 73726 86658
rect 73726 86606 73778 86658
rect 73778 86606 73780 86658
rect 73724 86604 73780 86606
rect 73388 86098 73444 86100
rect 73388 86046 73390 86098
rect 73390 86046 73442 86098
rect 73442 86046 73444 86098
rect 73388 86044 73444 86046
rect 74396 86658 74452 86660
rect 74396 86606 74398 86658
rect 74398 86606 74450 86658
rect 74450 86606 74452 86658
rect 74396 86604 74452 86606
rect 73164 85596 73220 85652
rect 73948 84476 74004 84532
rect 73612 84306 73668 84308
rect 73612 84254 73614 84306
rect 73614 84254 73666 84306
rect 73666 84254 73668 84306
rect 73612 84252 73668 84254
rect 74620 84252 74676 84308
rect 74732 85708 74788 85764
rect 75516 86604 75572 86660
rect 74956 86492 75012 86548
rect 75292 85708 75348 85764
rect 75740 86546 75796 86548
rect 75740 86494 75742 86546
rect 75742 86494 75794 86546
rect 75794 86494 75796 86546
rect 75740 86492 75796 86494
rect 76524 85820 76580 85876
rect 74844 84924 74900 84980
rect 75628 84978 75684 84980
rect 75628 84926 75630 84978
rect 75630 84926 75682 84978
rect 75682 84926 75684 84978
rect 75628 84924 75684 84926
rect 75516 84252 75572 84308
rect 73164 83244 73220 83300
rect 73276 82572 73332 82628
rect 72828 81842 72884 81844
rect 72828 81790 72830 81842
rect 72830 81790 72882 81842
rect 72882 81790 72884 81842
rect 72828 81788 72884 81790
rect 75404 84028 75460 84084
rect 73836 82626 73892 82628
rect 73836 82574 73838 82626
rect 73838 82574 73890 82626
rect 73890 82574 73892 82626
rect 73836 82572 73892 82574
rect 74956 82572 75012 82628
rect 75404 82066 75460 82068
rect 75404 82014 75406 82066
rect 75406 82014 75458 82066
rect 75458 82014 75460 82066
rect 75404 82012 75460 82014
rect 73612 81788 73668 81844
rect 73276 81676 73332 81732
rect 73836 81730 73892 81732
rect 73836 81678 73838 81730
rect 73838 81678 73890 81730
rect 73890 81678 73892 81730
rect 73836 81676 73892 81678
rect 74284 81730 74340 81732
rect 74284 81678 74286 81730
rect 74286 81678 74338 81730
rect 74338 81678 74340 81730
rect 74284 81676 74340 81678
rect 74844 81730 74900 81732
rect 74844 81678 74846 81730
rect 74846 81678 74898 81730
rect 74898 81678 74900 81730
rect 74844 81676 74900 81678
rect 73836 81394 73892 81396
rect 73836 81342 73838 81394
rect 73838 81342 73890 81394
rect 73890 81342 73892 81394
rect 73836 81340 73892 81342
rect 71708 80892 71764 80948
rect 71708 80108 71764 80164
rect 72268 79826 72324 79828
rect 72268 79774 72270 79826
rect 72270 79774 72322 79826
rect 72322 79774 72324 79826
rect 72268 79772 72324 79774
rect 71708 78652 71764 78708
rect 70812 77250 70868 77252
rect 70812 77198 70814 77250
rect 70814 77198 70866 77250
rect 70866 77198 70868 77250
rect 70812 77196 70868 77198
rect 70588 76412 70644 76468
rect 69692 75068 69748 75124
rect 70588 75122 70644 75124
rect 70588 75070 70590 75122
rect 70590 75070 70642 75122
rect 70642 75070 70644 75122
rect 70588 75068 70644 75070
rect 71820 77250 71876 77252
rect 71820 77198 71822 77250
rect 71822 77198 71874 77250
rect 71874 77198 71876 77250
rect 71820 77196 71876 77198
rect 71260 76412 71316 76468
rect 71260 75794 71316 75796
rect 71260 75742 71262 75794
rect 71262 75742 71314 75794
rect 71314 75742 71316 75794
rect 71260 75740 71316 75742
rect 71932 76300 71988 76356
rect 71596 75740 71652 75796
rect 72604 77868 72660 77924
rect 73836 80108 73892 80164
rect 76076 85708 76132 85764
rect 77868 86044 77924 86100
rect 77420 85762 77476 85764
rect 77420 85710 77422 85762
rect 77422 85710 77474 85762
rect 77474 85710 77476 85762
rect 77420 85708 77476 85710
rect 78204 85708 78260 85764
rect 77420 84306 77476 84308
rect 77420 84254 77422 84306
rect 77422 84254 77474 84306
rect 77474 84254 77476 84306
rect 77420 84252 77476 84254
rect 76412 84028 76468 84084
rect 77420 84028 77476 84084
rect 76412 83410 76468 83412
rect 76412 83358 76414 83410
rect 76414 83358 76466 83410
rect 76466 83358 76468 83410
rect 76412 83356 76468 83358
rect 77532 82236 77588 82292
rect 77532 82012 77588 82068
rect 77868 82066 77924 82068
rect 77868 82014 77870 82066
rect 77870 82014 77922 82066
rect 77922 82014 77924 82066
rect 77868 82012 77924 82014
rect 75740 81676 75796 81732
rect 76524 81730 76580 81732
rect 76524 81678 76526 81730
rect 76526 81678 76578 81730
rect 76578 81678 76580 81730
rect 76524 81676 76580 81678
rect 77196 81676 77252 81732
rect 75068 81394 75124 81396
rect 75068 81342 75070 81394
rect 75070 81342 75122 81394
rect 75122 81342 75124 81394
rect 75068 81340 75124 81342
rect 75292 81340 75348 81396
rect 74732 80668 74788 80724
rect 74508 80498 74564 80500
rect 74508 80446 74510 80498
rect 74510 80446 74562 80498
rect 74562 80446 74564 80498
rect 74508 80444 74564 80446
rect 74172 78652 74228 78708
rect 73164 77868 73220 77924
rect 72940 77756 72996 77812
rect 72156 77138 72212 77140
rect 72156 77086 72158 77138
rect 72158 77086 72210 77138
rect 72210 77086 72212 77138
rect 72156 77084 72212 77086
rect 72716 77138 72772 77140
rect 72716 77086 72718 77138
rect 72718 77086 72770 77138
rect 72770 77086 72772 77138
rect 72716 77084 72772 77086
rect 72156 76860 72212 76916
rect 72604 76354 72660 76356
rect 72604 76302 72606 76354
rect 72606 76302 72658 76354
rect 72658 76302 72660 76354
rect 72604 76300 72660 76302
rect 72156 76076 72212 76132
rect 72828 76188 72884 76244
rect 72044 75740 72100 75796
rect 71932 75628 71988 75684
rect 70588 74002 70644 74004
rect 70588 73950 70590 74002
rect 70590 73950 70642 74002
rect 70642 73950 70644 74002
rect 70588 73948 70644 73950
rect 70028 73836 70084 73892
rect 71260 73890 71316 73892
rect 71260 73838 71262 73890
rect 71262 73838 71314 73890
rect 71314 73838 71316 73890
rect 71260 73836 71316 73838
rect 69804 73164 69860 73220
rect 71148 73218 71204 73220
rect 71148 73166 71150 73218
rect 71150 73166 71202 73218
rect 71202 73166 71204 73218
rect 71148 73164 71204 73166
rect 70812 72434 70868 72436
rect 70812 72382 70814 72434
rect 70814 72382 70866 72434
rect 70866 72382 70868 72434
rect 70812 72380 70868 72382
rect 68572 70866 68628 70868
rect 68572 70814 68574 70866
rect 68574 70814 68626 70866
rect 68626 70814 68628 70866
rect 68572 70812 68628 70814
rect 68684 69580 68740 69636
rect 68796 70700 68852 70756
rect 68348 68236 68404 68292
rect 68460 67730 68516 67732
rect 68460 67678 68462 67730
rect 68462 67678 68514 67730
rect 68514 67678 68516 67730
rect 68460 67676 68516 67678
rect 67564 67564 67620 67620
rect 68572 67452 68628 67508
rect 68684 67340 68740 67396
rect 69580 71036 69636 71092
rect 69132 70476 69188 70532
rect 69244 69522 69300 69524
rect 69244 69470 69246 69522
rect 69246 69470 69298 69522
rect 69298 69470 69300 69522
rect 69244 69468 69300 69470
rect 71036 70082 71092 70084
rect 71036 70030 71038 70082
rect 71038 70030 71090 70082
rect 71090 70030 71092 70082
rect 71036 70028 71092 70030
rect 70252 69634 70308 69636
rect 70252 69582 70254 69634
rect 70254 69582 70306 69634
rect 70306 69582 70308 69634
rect 70252 69580 70308 69582
rect 69356 69356 69412 69412
rect 70588 68796 70644 68852
rect 69916 68514 69972 68516
rect 69916 68462 69918 68514
rect 69918 68462 69970 68514
rect 69970 68462 69972 68514
rect 69916 68460 69972 68462
rect 69580 68348 69636 68404
rect 69020 67676 69076 67732
rect 67452 66892 67508 66948
rect 67340 64876 67396 64932
rect 67340 64652 67396 64708
rect 67340 64316 67396 64372
rect 67340 63868 67396 63924
rect 67788 66780 67844 66836
rect 68572 66274 68628 66276
rect 68572 66222 68574 66274
rect 68574 66222 68626 66274
rect 68626 66222 68628 66274
rect 68572 66220 68628 66222
rect 67900 66162 67956 66164
rect 67900 66110 67902 66162
rect 67902 66110 67954 66162
rect 67954 66110 67956 66162
rect 67900 66108 67956 66110
rect 67788 65100 67844 65156
rect 67676 64652 67732 64708
rect 68348 65324 68404 65380
rect 68124 64876 68180 64932
rect 68236 64540 68292 64596
rect 68348 63922 68404 63924
rect 68348 63870 68350 63922
rect 68350 63870 68402 63922
rect 68402 63870 68404 63922
rect 68348 63868 68404 63870
rect 68460 64876 68516 64932
rect 68572 64594 68628 64596
rect 68572 64542 68574 64594
rect 68574 64542 68626 64594
rect 68626 64542 68628 64594
rect 68572 64540 68628 64542
rect 68796 66780 68852 66836
rect 70588 68236 70644 68292
rect 69580 67452 69636 67508
rect 69468 66946 69524 66948
rect 69468 66894 69470 66946
rect 69470 66894 69522 66946
rect 69522 66894 69524 66946
rect 69468 66892 69524 66894
rect 69916 67340 69972 67396
rect 70252 67170 70308 67172
rect 70252 67118 70254 67170
rect 70254 67118 70306 67170
rect 70306 67118 70308 67170
rect 70252 67116 70308 67118
rect 70140 66892 70196 66948
rect 69804 66220 69860 66276
rect 69692 66162 69748 66164
rect 69692 66110 69694 66162
rect 69694 66110 69746 66162
rect 69746 66110 69748 66162
rect 69692 66108 69748 66110
rect 69468 65884 69524 65940
rect 69804 65884 69860 65940
rect 69244 65660 69300 65716
rect 69692 65100 69748 65156
rect 70364 64988 70420 65044
rect 69356 64594 69412 64596
rect 69356 64542 69358 64594
rect 69358 64542 69410 64594
rect 69410 64542 69412 64594
rect 69356 64540 69412 64542
rect 68908 64204 68964 64260
rect 69244 63026 69300 63028
rect 69244 62974 69246 63026
rect 69246 62974 69298 63026
rect 69298 62974 69300 63026
rect 69244 62972 69300 62974
rect 68908 62748 68964 62804
rect 70476 64876 70532 64932
rect 70700 67116 70756 67172
rect 71708 74620 71764 74676
rect 71484 73948 71540 74004
rect 72268 74620 72324 74676
rect 72268 74002 72324 74004
rect 72268 73950 72270 74002
rect 72270 73950 72322 74002
rect 72322 73950 72324 74002
rect 72268 73948 72324 73950
rect 72716 74002 72772 74004
rect 72716 73950 72718 74002
rect 72718 73950 72770 74002
rect 72770 73950 72772 74002
rect 72716 73948 72772 73950
rect 71708 73836 71764 73892
rect 72156 72380 72212 72436
rect 72044 71596 72100 71652
rect 71372 71090 71428 71092
rect 71372 71038 71374 71090
rect 71374 71038 71426 71090
rect 71426 71038 71428 71090
rect 71372 71036 71428 71038
rect 71484 70812 71540 70868
rect 71372 70588 71428 70644
rect 72044 70588 72100 70644
rect 71484 69580 71540 69636
rect 72268 72044 72324 72100
rect 72604 71932 72660 71988
rect 71372 69298 71428 69300
rect 71372 69246 71374 69298
rect 71374 69246 71426 69298
rect 71426 69246 71428 69298
rect 71372 69244 71428 69246
rect 72828 70028 72884 70084
rect 72492 69634 72548 69636
rect 72492 69582 72494 69634
rect 72494 69582 72546 69634
rect 72546 69582 72548 69634
rect 72492 69580 72548 69582
rect 72380 69244 72436 69300
rect 71372 68124 71428 68180
rect 71820 68460 71876 68516
rect 71148 66780 71204 66836
rect 70700 65548 70756 65604
rect 70812 66108 70868 66164
rect 71036 65996 71092 66052
rect 70924 65772 70980 65828
rect 71148 65490 71204 65492
rect 71148 65438 71150 65490
rect 71150 65438 71202 65490
rect 71202 65438 71204 65490
rect 71148 65436 71204 65438
rect 71596 67618 71652 67620
rect 71596 67566 71598 67618
rect 71598 67566 71650 67618
rect 71650 67566 71652 67618
rect 71596 67564 71652 67566
rect 72492 68236 72548 68292
rect 73052 69298 73108 69300
rect 73052 69246 73054 69298
rect 73054 69246 73106 69298
rect 73106 69246 73108 69298
rect 73052 69244 73108 69246
rect 72044 67618 72100 67620
rect 72044 67566 72046 67618
rect 72046 67566 72098 67618
rect 72098 67566 72100 67618
rect 72044 67564 72100 67566
rect 72268 67564 72324 67620
rect 72156 66892 72212 66948
rect 71932 66668 71988 66724
rect 72044 65378 72100 65380
rect 72044 65326 72046 65378
rect 72046 65326 72098 65378
rect 72098 65326 72100 65378
rect 72044 65324 72100 65326
rect 71260 64876 71316 64932
rect 70588 64034 70644 64036
rect 70588 63982 70590 64034
rect 70590 63982 70642 64034
rect 70642 63982 70644 64034
rect 70588 63980 70644 63982
rect 70700 63644 70756 63700
rect 69916 62972 69972 63028
rect 68236 61628 68292 61684
rect 67452 61570 67508 61572
rect 67452 61518 67454 61570
rect 67454 61518 67506 61570
rect 67506 61518 67508 61570
rect 67452 61516 67508 61518
rect 67676 61458 67732 61460
rect 67676 61406 67678 61458
rect 67678 61406 67730 61458
rect 67730 61406 67732 61458
rect 67676 61404 67732 61406
rect 67116 60732 67172 60788
rect 66780 59890 66836 59892
rect 66780 59838 66782 59890
rect 66782 59838 66834 59890
rect 66834 59838 66836 59890
rect 66780 59836 66836 59838
rect 65772 59052 65828 59108
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65884 58380 65940 58436
rect 65660 58156 65716 58212
rect 66108 58156 66164 58212
rect 65548 57874 65604 57876
rect 65548 57822 65550 57874
rect 65550 57822 65602 57874
rect 65602 57822 65604 57874
rect 65548 57820 65604 57822
rect 66444 58210 66500 58212
rect 66444 58158 66446 58210
rect 66446 58158 66498 58210
rect 66498 58158 66500 58210
rect 66444 58156 66500 58158
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 64764 57036 64820 57092
rect 65548 56194 65604 56196
rect 65548 56142 65550 56194
rect 65550 56142 65602 56194
rect 65602 56142 65604 56194
rect 65548 56140 65604 56142
rect 64764 55132 64820 55188
rect 66444 55804 66500 55860
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 65324 55020 65380 55076
rect 65324 54684 65380 54740
rect 65660 55132 65716 55188
rect 66892 59052 66948 59108
rect 67004 58492 67060 58548
rect 66892 58210 66948 58212
rect 66892 58158 66894 58210
rect 66894 58158 66946 58210
rect 66946 58158 66948 58210
rect 66892 58156 66948 58158
rect 66892 56700 66948 56756
rect 67228 60114 67284 60116
rect 67228 60062 67230 60114
rect 67230 60062 67282 60114
rect 67282 60062 67284 60114
rect 67228 60060 67284 60062
rect 67564 60396 67620 60452
rect 67676 60732 67732 60788
rect 67340 59948 67396 60004
rect 68012 60508 68068 60564
rect 67116 56588 67172 56644
rect 68460 61682 68516 61684
rect 68460 61630 68462 61682
rect 68462 61630 68514 61682
rect 68514 61630 68516 61682
rect 68460 61628 68516 61630
rect 69244 61740 69300 61796
rect 69244 61404 69300 61460
rect 68460 60396 68516 60452
rect 68572 59948 68628 60004
rect 68572 59724 68628 59780
rect 68460 59500 68516 59556
rect 68124 58492 68180 58548
rect 68236 58434 68292 58436
rect 68236 58382 68238 58434
rect 68238 58382 68290 58434
rect 68290 58382 68292 58434
rect 68236 58380 68292 58382
rect 68124 57484 68180 57540
rect 65548 53788 65604 53844
rect 64540 53564 64596 53620
rect 65660 53618 65716 53620
rect 65660 53566 65662 53618
rect 65662 53566 65714 53618
rect 65714 53566 65716 53618
rect 65660 53564 65716 53566
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 66108 53618 66164 53620
rect 66108 53566 66110 53618
rect 66110 53566 66162 53618
rect 66162 53566 66164 53618
rect 66108 53564 66164 53566
rect 64540 53058 64596 53060
rect 64540 53006 64542 53058
rect 64542 53006 64594 53058
rect 64594 53006 64596 53058
rect 64540 53004 64596 53006
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 64764 51548 64820 51604
rect 64540 51324 64596 51380
rect 65324 51602 65380 51604
rect 65324 51550 65326 51602
rect 65326 51550 65378 51602
rect 65378 51550 65380 51602
rect 65324 51548 65380 51550
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 64540 50428 64596 50484
rect 65324 50482 65380 50484
rect 65324 50430 65326 50482
rect 65326 50430 65378 50482
rect 65378 50430 65380 50482
rect 65324 50428 65380 50430
rect 65436 50370 65492 50372
rect 65436 50318 65438 50370
rect 65438 50318 65490 50370
rect 65490 50318 65492 50370
rect 65436 50316 65492 50318
rect 65324 49810 65380 49812
rect 65324 49758 65326 49810
rect 65326 49758 65378 49810
rect 65378 49758 65380 49810
rect 65324 49756 65380 49758
rect 64652 49698 64708 49700
rect 64652 49646 64654 49698
rect 64654 49646 64706 49698
rect 64706 49646 64708 49698
rect 64652 49644 64708 49646
rect 65436 49644 65492 49700
rect 65996 50316 66052 50372
rect 66444 50428 66500 50484
rect 67004 53730 67060 53732
rect 67004 53678 67006 53730
rect 67006 53678 67058 53730
rect 67058 53678 67060 53730
rect 67004 53676 67060 53678
rect 67452 55858 67508 55860
rect 67452 55806 67454 55858
rect 67454 55806 67506 55858
rect 67506 55806 67508 55858
rect 67452 55804 67508 55806
rect 68572 59276 68628 59332
rect 68572 58434 68628 58436
rect 68572 58382 68574 58434
rect 68574 58382 68626 58434
rect 68626 58382 68628 58434
rect 68572 58380 68628 58382
rect 68348 56082 68404 56084
rect 68348 56030 68350 56082
rect 68350 56030 68402 56082
rect 68402 56030 68404 56082
rect 68348 56028 68404 56030
rect 68124 55356 68180 55412
rect 68572 55692 68628 55748
rect 67788 53730 67844 53732
rect 67788 53678 67790 53730
rect 67790 53678 67842 53730
rect 67842 53678 67844 53730
rect 67788 53676 67844 53678
rect 67340 53058 67396 53060
rect 67340 53006 67342 53058
rect 67342 53006 67394 53058
rect 67394 53006 67396 53058
rect 67340 53004 67396 53006
rect 67004 52556 67060 52612
rect 67116 52444 67172 52500
rect 68236 53004 68292 53060
rect 68572 53452 68628 53508
rect 68572 52444 68628 52500
rect 67788 52050 67844 52052
rect 67788 51998 67790 52050
rect 67790 51998 67842 52050
rect 67842 51998 67844 52050
rect 67788 51996 67844 51998
rect 68572 52108 68628 52164
rect 67340 50540 67396 50596
rect 66332 49922 66388 49924
rect 66332 49870 66334 49922
rect 66334 49870 66386 49922
rect 66386 49870 66388 49922
rect 66332 49868 66388 49870
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65212 48914 65268 48916
rect 65212 48862 65214 48914
rect 65214 48862 65266 48914
rect 65266 48862 65268 48914
rect 65212 48860 65268 48862
rect 65100 48524 65156 48580
rect 64876 47180 64932 47236
rect 65548 48354 65604 48356
rect 65548 48302 65550 48354
rect 65550 48302 65602 48354
rect 65602 48302 65604 48354
rect 65548 48300 65604 48302
rect 65436 48076 65492 48132
rect 66444 49532 66500 49588
rect 66892 49922 66948 49924
rect 66892 49870 66894 49922
rect 66894 49870 66946 49922
rect 66946 49870 66948 49922
rect 66892 49868 66948 49870
rect 66892 48636 66948 48692
rect 66332 48524 66388 48580
rect 68572 50540 68628 50596
rect 68236 49868 68292 49924
rect 68012 49810 68068 49812
rect 68012 49758 68014 49810
rect 68014 49758 68066 49810
rect 68066 49758 68068 49810
rect 68012 49756 68068 49758
rect 67452 49532 67508 49588
rect 67228 48972 67284 49028
rect 65884 48188 65940 48244
rect 66108 48242 66164 48244
rect 66108 48190 66110 48242
rect 66110 48190 66162 48242
rect 66162 48190 66164 48242
rect 66108 48188 66164 48190
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 66108 47404 66164 47460
rect 65660 47180 65716 47236
rect 66220 47234 66276 47236
rect 66220 47182 66222 47234
rect 66222 47182 66274 47234
rect 66274 47182 66276 47234
rect 66220 47180 66276 47182
rect 67116 48412 67172 48468
rect 66556 47458 66612 47460
rect 66556 47406 66558 47458
rect 66558 47406 66610 47458
rect 66610 47406 66612 47458
rect 66556 47404 66612 47406
rect 66332 47068 66388 47124
rect 65548 46786 65604 46788
rect 65548 46734 65550 46786
rect 65550 46734 65602 46786
rect 65602 46734 65604 46786
rect 65548 46732 65604 46734
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65324 45388 65380 45444
rect 66444 44940 66500 44996
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 64204 43596 64260 43652
rect 64540 43538 64596 43540
rect 64540 43486 64542 43538
rect 64542 43486 64594 43538
rect 64594 43486 64596 43538
rect 64540 43484 64596 43486
rect 64428 43260 64484 43316
rect 63868 42866 63924 42868
rect 63868 42814 63870 42866
rect 63870 42814 63922 42866
rect 63922 42814 63924 42866
rect 63868 42812 63924 42814
rect 63420 41858 63476 41860
rect 63420 41806 63422 41858
rect 63422 41806 63474 41858
rect 63474 41806 63476 41858
rect 63420 41804 63476 41806
rect 63532 40514 63588 40516
rect 63532 40462 63534 40514
rect 63534 40462 63586 40514
rect 63586 40462 63588 40514
rect 63532 40460 63588 40462
rect 64316 41692 64372 41748
rect 64204 41244 64260 41300
rect 63980 40514 64036 40516
rect 63980 40462 63982 40514
rect 63982 40462 64034 40514
rect 64034 40462 64036 40514
rect 63980 40460 64036 40462
rect 64316 41468 64372 41524
rect 64428 41244 64484 41300
rect 64652 41804 64708 41860
rect 63756 39340 63812 39396
rect 63980 38946 64036 38948
rect 63980 38894 63982 38946
rect 63982 38894 64034 38946
rect 64034 38894 64036 38946
rect 63980 38892 64036 38894
rect 63420 38780 63476 38836
rect 64204 38834 64260 38836
rect 64204 38782 64206 38834
rect 64206 38782 64258 38834
rect 64258 38782 64260 38834
rect 64204 38780 64260 38782
rect 66332 43596 66388 43652
rect 65324 43484 65380 43540
rect 64988 41186 65044 41188
rect 64988 41134 64990 41186
rect 64990 41134 65042 41186
rect 65042 41134 65044 41186
rect 64988 41132 65044 41134
rect 65212 40460 65268 40516
rect 65772 43538 65828 43540
rect 65772 43486 65774 43538
rect 65774 43486 65826 43538
rect 65826 43486 65828 43538
rect 65772 43484 65828 43486
rect 65772 43260 65828 43316
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65772 42082 65828 42084
rect 65772 42030 65774 42082
rect 65774 42030 65826 42082
rect 65826 42030 65828 42082
rect 65772 42028 65828 42030
rect 66892 48130 66948 48132
rect 66892 48078 66894 48130
rect 66894 48078 66946 48130
rect 66946 48078 66948 48130
rect 66892 48076 66948 48078
rect 66892 47852 66948 47908
rect 67004 47404 67060 47460
rect 67004 45106 67060 45108
rect 67004 45054 67006 45106
rect 67006 45054 67058 45106
rect 67058 45054 67060 45106
rect 67004 45052 67060 45054
rect 66780 43484 66836 43540
rect 67452 48860 67508 48916
rect 67340 48466 67396 48468
rect 67340 48414 67342 48466
rect 67342 48414 67394 48466
rect 67394 48414 67396 48466
rect 67340 48412 67396 48414
rect 67452 48076 67508 48132
rect 68236 48860 68292 48916
rect 70140 62354 70196 62356
rect 70140 62302 70142 62354
rect 70142 62302 70194 62354
rect 70194 62302 70196 62354
rect 70140 62300 70196 62302
rect 69916 62188 69972 62244
rect 69692 61516 69748 61572
rect 70252 61570 70308 61572
rect 70252 61518 70254 61570
rect 70254 61518 70306 61570
rect 70306 61518 70308 61570
rect 70252 61516 70308 61518
rect 70028 61180 70084 61236
rect 69916 60844 69972 60900
rect 69356 60786 69412 60788
rect 69356 60734 69358 60786
rect 69358 60734 69410 60786
rect 69410 60734 69412 60786
rect 69356 60732 69412 60734
rect 69244 60562 69300 60564
rect 69244 60510 69246 60562
rect 69246 60510 69298 60562
rect 69298 60510 69300 60562
rect 69244 60508 69300 60510
rect 69804 60396 69860 60452
rect 69468 60002 69524 60004
rect 69468 59950 69470 60002
rect 69470 59950 69522 60002
rect 69522 59950 69524 60002
rect 69468 59948 69524 59950
rect 69356 59330 69412 59332
rect 69356 59278 69358 59330
rect 69358 59278 69410 59330
rect 69410 59278 69412 59330
rect 69356 59276 69412 59278
rect 69244 59052 69300 59108
rect 69244 58492 69300 58548
rect 68796 57538 68852 57540
rect 68796 57486 68798 57538
rect 68798 57486 68850 57538
rect 68850 57486 68852 57538
rect 68796 57484 68852 57486
rect 68908 56082 68964 56084
rect 68908 56030 68910 56082
rect 68910 56030 68962 56082
rect 68962 56030 68964 56082
rect 68908 56028 68964 56030
rect 71260 64706 71316 64708
rect 71260 64654 71262 64706
rect 71262 64654 71314 64706
rect 71314 64654 71316 64706
rect 71260 64652 71316 64654
rect 72044 64876 72100 64932
rect 71596 64706 71652 64708
rect 71596 64654 71598 64706
rect 71598 64654 71650 64706
rect 71650 64654 71652 64706
rect 71596 64652 71652 64654
rect 70476 62300 70532 62356
rect 70924 63644 70980 63700
rect 70476 61458 70532 61460
rect 70476 61406 70478 61458
rect 70478 61406 70530 61458
rect 70530 61406 70532 61458
rect 70476 61404 70532 61406
rect 71036 63532 71092 63588
rect 71036 62636 71092 62692
rect 71036 62354 71092 62356
rect 71036 62302 71038 62354
rect 71038 62302 71090 62354
rect 71090 62302 71092 62354
rect 71036 62300 71092 62302
rect 70924 62188 70980 62244
rect 70700 61180 70756 61236
rect 70140 60898 70196 60900
rect 70140 60846 70142 60898
rect 70142 60846 70194 60898
rect 70194 60846 70196 60898
rect 70140 60844 70196 60846
rect 71372 63644 71428 63700
rect 71148 62076 71204 62132
rect 71708 64092 71764 64148
rect 72492 66108 72548 66164
rect 72604 66050 72660 66052
rect 72604 65998 72606 66050
rect 72606 65998 72658 66050
rect 72658 65998 72660 66050
rect 72604 65996 72660 65998
rect 73052 65548 73108 65604
rect 72604 65436 72660 65492
rect 72044 63980 72100 64036
rect 71708 63868 71764 63924
rect 70028 60732 70084 60788
rect 71148 61570 71204 61572
rect 71148 61518 71150 61570
rect 71150 61518 71202 61570
rect 71202 61518 71204 61570
rect 71148 61516 71204 61518
rect 69916 60060 69972 60116
rect 69468 58268 69524 58324
rect 69580 58604 69636 58660
rect 69692 57148 69748 57204
rect 69356 56028 69412 56084
rect 70252 59724 70308 59780
rect 70700 60508 70756 60564
rect 70476 59724 70532 59780
rect 70588 59500 70644 59556
rect 70476 59052 70532 59108
rect 70252 58546 70308 58548
rect 70252 58494 70254 58546
rect 70254 58494 70306 58546
rect 70306 58494 70308 58546
rect 70252 58492 70308 58494
rect 70140 57932 70196 57988
rect 70364 57874 70420 57876
rect 70364 57822 70366 57874
rect 70366 57822 70418 57874
rect 70418 57822 70420 57874
rect 70364 57820 70420 57822
rect 70140 57148 70196 57204
rect 68684 49756 68740 49812
rect 69244 53506 69300 53508
rect 69244 53454 69246 53506
rect 69246 53454 69298 53506
rect 69298 53454 69300 53506
rect 69244 53452 69300 53454
rect 69132 52108 69188 52164
rect 68684 49196 68740 49252
rect 69468 54626 69524 54628
rect 69468 54574 69470 54626
rect 69470 54574 69522 54626
rect 69522 54574 69524 54626
rect 69468 54572 69524 54574
rect 69580 53340 69636 53396
rect 69916 54626 69972 54628
rect 69916 54574 69918 54626
rect 69918 54574 69970 54626
rect 69970 54574 69972 54626
rect 69916 54572 69972 54574
rect 70028 52556 70084 52612
rect 70364 53452 70420 53508
rect 70364 53170 70420 53172
rect 70364 53118 70366 53170
rect 70366 53118 70418 53170
rect 70418 53118 70420 53170
rect 70364 53116 70420 53118
rect 70140 52162 70196 52164
rect 70140 52110 70142 52162
rect 70142 52110 70194 52162
rect 70194 52110 70196 52162
rect 70140 52108 70196 52110
rect 70812 59948 70868 60004
rect 70812 58604 70868 58660
rect 70924 59500 70980 59556
rect 70588 57484 70644 57540
rect 70812 57538 70868 57540
rect 70812 57486 70814 57538
rect 70814 57486 70866 57538
rect 70866 57486 70868 57538
rect 70812 57484 70868 57486
rect 70588 56978 70644 56980
rect 70588 56926 70590 56978
rect 70590 56926 70642 56978
rect 70642 56926 70644 56978
rect 70588 56924 70644 56926
rect 71932 63922 71988 63924
rect 71932 63870 71934 63922
rect 71934 63870 71986 63922
rect 71986 63870 71988 63922
rect 71932 63868 71988 63870
rect 72380 64034 72436 64036
rect 72380 63982 72382 64034
rect 72382 63982 72434 64034
rect 72434 63982 72436 64034
rect 72380 63980 72436 63982
rect 72156 63868 72212 63924
rect 72268 63756 72324 63812
rect 71484 62242 71540 62244
rect 71484 62190 71486 62242
rect 71486 62190 71538 62242
rect 71538 62190 71540 62242
rect 71484 62188 71540 62190
rect 71372 60898 71428 60900
rect 71372 60846 71374 60898
rect 71374 60846 71426 60898
rect 71426 60846 71428 60898
rect 71372 60844 71428 60846
rect 71932 62636 71988 62692
rect 71708 62076 71764 62132
rect 72716 65378 72772 65380
rect 72716 65326 72718 65378
rect 72718 65326 72770 65378
rect 72770 65326 72772 65378
rect 72716 65324 72772 65326
rect 73948 77196 74004 77252
rect 73724 76188 73780 76244
rect 73388 75794 73444 75796
rect 73388 75742 73390 75794
rect 73390 75742 73442 75794
rect 73442 75742 73444 75794
rect 73388 75740 73444 75742
rect 73724 75628 73780 75684
rect 73724 74844 73780 74900
rect 73500 74620 73556 74676
rect 73276 73948 73332 74004
rect 73724 73948 73780 74004
rect 73836 72044 73892 72100
rect 73612 71932 73668 71988
rect 73276 71650 73332 71652
rect 73276 71598 73278 71650
rect 73278 71598 73330 71650
rect 73330 71598 73332 71650
rect 73276 71596 73332 71598
rect 73276 70924 73332 70980
rect 73836 71596 73892 71652
rect 74060 69244 74116 69300
rect 73500 68684 73556 68740
rect 73724 68684 73780 68740
rect 73388 68236 73444 68292
rect 73724 68236 73780 68292
rect 73388 67340 73444 67396
rect 73500 66892 73556 66948
rect 73276 65996 73332 66052
rect 73948 68124 74004 68180
rect 74060 69020 74116 69076
rect 73836 67842 73892 67844
rect 73836 67790 73838 67842
rect 73838 67790 73890 67842
rect 73890 67790 73892 67842
rect 73836 67788 73892 67790
rect 73948 67170 74004 67172
rect 73948 67118 73950 67170
rect 73950 67118 74002 67170
rect 74002 67118 74004 67170
rect 73948 67116 74004 67118
rect 74060 66274 74116 66276
rect 74060 66222 74062 66274
rect 74062 66222 74114 66274
rect 74114 66222 74116 66274
rect 74060 66220 74116 66222
rect 73724 66162 73780 66164
rect 73724 66110 73726 66162
rect 73726 66110 73778 66162
rect 73778 66110 73780 66162
rect 73724 66108 73780 66110
rect 73612 65996 73668 66052
rect 73948 65436 74004 65492
rect 72604 63756 72660 63812
rect 72716 63868 72772 63924
rect 72380 61852 72436 61908
rect 72492 61964 72548 62020
rect 71484 60508 71540 60564
rect 72268 61570 72324 61572
rect 72268 61518 72270 61570
rect 72270 61518 72322 61570
rect 72322 61518 72324 61570
rect 72268 61516 72324 61518
rect 71932 60002 71988 60004
rect 71932 59950 71934 60002
rect 71934 59950 71986 60002
rect 71986 59950 71988 60002
rect 71932 59948 71988 59950
rect 72156 60844 72212 60900
rect 71484 59276 71540 59332
rect 70924 56364 70980 56420
rect 70700 54572 70756 54628
rect 70924 53452 70980 53508
rect 70812 53340 70868 53396
rect 70812 52332 70868 52388
rect 70700 51996 70756 52052
rect 71372 58716 71428 58772
rect 71484 58604 71540 58660
rect 72156 60508 72212 60564
rect 71596 58268 71652 58324
rect 71820 58322 71876 58324
rect 71820 58270 71822 58322
rect 71822 58270 71874 58322
rect 71874 58270 71876 58322
rect 71820 58268 71876 58270
rect 72268 60284 72324 60340
rect 72044 58716 72100 58772
rect 71820 58044 71876 58100
rect 71372 57484 71428 57540
rect 71148 57036 71204 57092
rect 71148 56642 71204 56644
rect 71148 56590 71150 56642
rect 71150 56590 71202 56642
rect 71202 56590 71204 56642
rect 71148 56588 71204 56590
rect 71484 56476 71540 56532
rect 72156 58156 72212 58212
rect 72044 56476 72100 56532
rect 71932 56306 71988 56308
rect 71932 56254 71934 56306
rect 71934 56254 71986 56306
rect 71986 56254 71988 56306
rect 71932 56252 71988 56254
rect 71148 54626 71204 54628
rect 71148 54574 71150 54626
rect 71150 54574 71202 54626
rect 71202 54574 71204 54626
rect 71148 54572 71204 54574
rect 72492 60844 72548 60900
rect 72828 61852 72884 61908
rect 72828 61458 72884 61460
rect 72828 61406 72830 61458
rect 72830 61406 72882 61458
rect 72882 61406 72884 61458
rect 72828 61404 72884 61406
rect 73276 61852 73332 61908
rect 72940 61180 72996 61236
rect 72716 60284 72772 60340
rect 72604 59948 72660 60004
rect 73724 65324 73780 65380
rect 74060 64652 74116 64708
rect 74956 77756 75012 77812
rect 74732 77084 74788 77140
rect 74284 77026 74340 77028
rect 74284 76974 74286 77026
rect 74286 76974 74338 77026
rect 74338 76974 74340 77026
rect 74284 76972 74340 76974
rect 74284 76188 74340 76244
rect 74396 76300 74452 76356
rect 74284 75740 74340 75796
rect 75180 80444 75236 80500
rect 75964 80556 76020 80612
rect 75180 78706 75236 78708
rect 75180 78654 75182 78706
rect 75182 78654 75234 78706
rect 75234 78654 75236 78706
rect 75180 78652 75236 78654
rect 74956 75628 75012 75684
rect 75068 75570 75124 75572
rect 75068 75518 75070 75570
rect 75070 75518 75122 75570
rect 75122 75518 75124 75570
rect 75068 75516 75124 75518
rect 74620 75122 74676 75124
rect 74620 75070 74622 75122
rect 74622 75070 74674 75122
rect 74674 75070 74676 75122
rect 74620 75068 74676 75070
rect 74396 74956 74452 75012
rect 75068 75010 75124 75012
rect 75068 74958 75070 75010
rect 75070 74958 75122 75010
rect 75122 74958 75124 75010
rect 75068 74956 75124 74958
rect 74284 74898 74340 74900
rect 74284 74846 74286 74898
rect 74286 74846 74338 74898
rect 74338 74846 74340 74898
rect 74284 74844 74340 74846
rect 74396 72156 74452 72212
rect 74284 71148 74340 71204
rect 75740 78764 75796 78820
rect 76188 80162 76244 80164
rect 76188 80110 76190 80162
rect 76190 80110 76242 80162
rect 76242 80110 76244 80162
rect 76188 80108 76244 80110
rect 78316 80668 78372 80724
rect 75516 78706 75572 78708
rect 75516 78654 75518 78706
rect 75518 78654 75570 78706
rect 75570 78654 75572 78706
rect 75516 78652 75572 78654
rect 76300 78706 76356 78708
rect 76300 78654 76302 78706
rect 76302 78654 76354 78706
rect 76354 78654 76356 78706
rect 76300 78652 76356 78654
rect 76748 78652 76804 78708
rect 77196 79490 77252 79492
rect 77196 79438 77198 79490
rect 77198 79438 77250 79490
rect 77250 79438 77252 79490
rect 77196 79436 77252 79438
rect 76188 78092 76244 78148
rect 76748 77980 76804 78036
rect 76524 77250 76580 77252
rect 76524 77198 76526 77250
rect 76526 77198 76578 77250
rect 76578 77198 76580 77250
rect 76524 77196 76580 77198
rect 76972 77196 77028 77252
rect 75516 76972 75572 77028
rect 75852 76636 75908 76692
rect 75404 76524 75460 76580
rect 75404 75740 75460 75796
rect 75964 75570 76020 75572
rect 75964 75518 75966 75570
rect 75966 75518 76018 75570
rect 76018 75518 76020 75570
rect 75964 75516 76020 75518
rect 76300 75682 76356 75684
rect 76300 75630 76302 75682
rect 76302 75630 76354 75682
rect 76354 75630 76356 75682
rect 76300 75628 76356 75630
rect 75964 75068 76020 75124
rect 75964 73164 76020 73220
rect 75180 72268 75236 72324
rect 75628 72044 75684 72100
rect 74844 71932 74900 71988
rect 75068 71596 75124 71652
rect 74956 69356 75012 69412
rect 74844 69298 74900 69300
rect 74844 69246 74846 69298
rect 74846 69246 74898 69298
rect 74898 69246 74900 69298
rect 74844 69244 74900 69246
rect 74732 69020 74788 69076
rect 74284 68796 74340 68852
rect 74284 68626 74340 68628
rect 74284 68574 74286 68626
rect 74286 68574 74338 68626
rect 74338 68574 74340 68626
rect 74284 68572 74340 68574
rect 74844 68348 74900 68404
rect 75628 71148 75684 71204
rect 75180 69804 75236 69860
rect 75516 70252 75572 70308
rect 81276 89402 81332 89404
rect 81276 89350 81278 89402
rect 81278 89350 81330 89402
rect 81330 89350 81332 89402
rect 81276 89348 81332 89350
rect 81380 89402 81436 89404
rect 81380 89350 81382 89402
rect 81382 89350 81434 89402
rect 81434 89350 81436 89402
rect 81380 89348 81436 89350
rect 81484 89402 81540 89404
rect 81484 89350 81486 89402
rect 81486 89350 81538 89402
rect 81538 89350 81540 89402
rect 81484 89348 81540 89350
rect 81276 87834 81332 87836
rect 81276 87782 81278 87834
rect 81278 87782 81330 87834
rect 81330 87782 81332 87834
rect 81276 87780 81332 87782
rect 81380 87834 81436 87836
rect 81380 87782 81382 87834
rect 81382 87782 81434 87834
rect 81434 87782 81436 87834
rect 81380 87780 81436 87782
rect 81484 87834 81540 87836
rect 81484 87782 81486 87834
rect 81486 87782 81538 87834
rect 81538 87782 81540 87834
rect 81484 87780 81540 87782
rect 79212 86098 79268 86100
rect 79212 86046 79214 86098
rect 79214 86046 79266 86098
rect 79266 86046 79268 86098
rect 79212 86044 79268 86046
rect 78540 83410 78596 83412
rect 78540 83358 78542 83410
rect 78542 83358 78594 83410
rect 78594 83358 78596 83410
rect 78540 83356 78596 83358
rect 78876 85762 78932 85764
rect 78876 85710 78878 85762
rect 78878 85710 78930 85762
rect 78930 85710 78932 85762
rect 78876 85708 78932 85710
rect 81228 86434 81284 86436
rect 81228 86382 81230 86434
rect 81230 86382 81282 86434
rect 81282 86382 81284 86434
rect 81228 86380 81284 86382
rect 81276 86266 81332 86268
rect 81276 86214 81278 86266
rect 81278 86214 81330 86266
rect 81330 86214 81332 86266
rect 81276 86212 81332 86214
rect 81380 86266 81436 86268
rect 81380 86214 81382 86266
rect 81382 86214 81434 86266
rect 81434 86214 81436 86266
rect 81380 86212 81436 86214
rect 81484 86266 81540 86268
rect 81484 86214 81486 86266
rect 81486 86214 81538 86266
rect 81538 86214 81540 86266
rect 81484 86212 81540 86214
rect 81900 86380 81956 86436
rect 79660 85708 79716 85764
rect 78764 84252 78820 84308
rect 79548 84252 79604 84308
rect 79772 85596 79828 85652
rect 80444 85596 80500 85652
rect 81676 85596 81732 85652
rect 81276 84698 81332 84700
rect 81276 84646 81278 84698
rect 81278 84646 81330 84698
rect 81330 84646 81332 84698
rect 81276 84644 81332 84646
rect 81380 84698 81436 84700
rect 81380 84646 81382 84698
rect 81382 84646 81434 84698
rect 81434 84646 81436 84698
rect 81380 84644 81436 84646
rect 81484 84698 81540 84700
rect 81484 84646 81486 84698
rect 81486 84646 81538 84698
rect 81538 84646 81540 84698
rect 81484 84644 81540 84646
rect 81676 84364 81732 84420
rect 80444 84252 80500 84308
rect 81452 84306 81508 84308
rect 81452 84254 81454 84306
rect 81454 84254 81506 84306
rect 81506 84254 81508 84306
rect 81452 84252 81508 84254
rect 80556 84140 80612 84196
rect 80444 83356 80500 83412
rect 79212 82236 79268 82292
rect 78652 82012 78708 82068
rect 80108 81170 80164 81172
rect 80108 81118 80110 81170
rect 80110 81118 80162 81170
rect 80162 81118 80164 81170
rect 80108 81116 80164 81118
rect 79548 80892 79604 80948
rect 79324 80668 79380 80724
rect 78876 79436 78932 79492
rect 78876 78988 78932 79044
rect 77308 78146 77364 78148
rect 77308 78094 77310 78146
rect 77310 78094 77362 78146
rect 77362 78094 77364 78146
rect 77308 78092 77364 78094
rect 77756 77308 77812 77364
rect 78092 78034 78148 78036
rect 78092 77982 78094 78034
rect 78094 77982 78146 78034
rect 78146 77982 78148 78034
rect 78092 77980 78148 77982
rect 77196 77138 77252 77140
rect 77196 77086 77198 77138
rect 77198 77086 77250 77138
rect 77250 77086 77252 77138
rect 77196 77084 77252 77086
rect 78316 77196 78372 77252
rect 77756 76690 77812 76692
rect 77756 76638 77758 76690
rect 77758 76638 77810 76690
rect 77810 76638 77812 76690
rect 77756 76636 77812 76638
rect 78316 76636 78372 76692
rect 77420 75628 77476 75684
rect 78540 77420 78596 77476
rect 78428 74844 78484 74900
rect 76524 73388 76580 73444
rect 76524 72044 76580 72100
rect 77196 73218 77252 73220
rect 77196 73166 77198 73218
rect 77198 73166 77250 73218
rect 77250 73166 77252 73218
rect 77196 73164 77252 73166
rect 77196 72322 77252 72324
rect 77196 72270 77198 72322
rect 77198 72270 77250 72322
rect 77250 72270 77252 72322
rect 77196 72268 77252 72270
rect 77868 73388 77924 73444
rect 78316 73164 78372 73220
rect 77420 72156 77476 72212
rect 76076 71596 76132 71652
rect 76076 70978 76132 70980
rect 76076 70926 76078 70978
rect 76078 70926 76130 70978
rect 76130 70926 76132 70978
rect 76076 70924 76132 70926
rect 76188 70306 76244 70308
rect 76188 70254 76190 70306
rect 76190 70254 76242 70306
rect 76242 70254 76244 70306
rect 76188 70252 76244 70254
rect 75740 69804 75796 69860
rect 76300 69468 76356 69524
rect 75404 69410 75460 69412
rect 75404 69358 75406 69410
rect 75406 69358 75458 69410
rect 75458 69358 75460 69410
rect 75404 69356 75460 69358
rect 75180 68796 75236 68852
rect 75740 68738 75796 68740
rect 75740 68686 75742 68738
rect 75742 68686 75794 68738
rect 75794 68686 75796 68738
rect 75740 68684 75796 68686
rect 74284 67676 74340 67732
rect 74508 67452 74564 67508
rect 74508 67282 74564 67284
rect 74508 67230 74510 67282
rect 74510 67230 74562 67282
rect 74562 67230 74564 67282
rect 74508 67228 74564 67230
rect 75068 67564 75124 67620
rect 74732 66892 74788 66948
rect 74732 66108 74788 66164
rect 74396 64706 74452 64708
rect 74396 64654 74398 64706
rect 74398 64654 74450 64706
rect 74450 64654 74452 64706
rect 74396 64652 74452 64654
rect 74060 62188 74116 62244
rect 73276 60508 73332 60564
rect 73500 60732 73556 60788
rect 72940 60226 72996 60228
rect 72940 60174 72942 60226
rect 72942 60174 72994 60226
rect 72994 60174 72996 60226
rect 72940 60172 72996 60174
rect 72828 58210 72884 58212
rect 72828 58158 72830 58210
rect 72830 58158 72882 58210
rect 72882 58158 72884 58210
rect 72828 58156 72884 58158
rect 72156 57036 72212 57092
rect 72156 56140 72212 56196
rect 72492 57596 72548 57652
rect 71148 53564 71204 53620
rect 71708 53564 71764 53620
rect 71260 53506 71316 53508
rect 71260 53454 71262 53506
rect 71262 53454 71314 53506
rect 71314 53454 71316 53506
rect 71260 53452 71316 53454
rect 72604 57538 72660 57540
rect 72604 57486 72606 57538
rect 72606 57486 72658 57538
rect 72658 57486 72660 57538
rect 72604 57484 72660 57486
rect 72604 56364 72660 56420
rect 72380 56194 72436 56196
rect 72380 56142 72382 56194
rect 72382 56142 72434 56194
rect 72434 56142 72436 56194
rect 72380 56140 72436 56142
rect 72268 54738 72324 54740
rect 72268 54686 72270 54738
rect 72270 54686 72322 54738
rect 72322 54686 72324 54738
rect 72268 54684 72324 54686
rect 72716 56252 72772 56308
rect 73052 58268 73108 58324
rect 73164 57820 73220 57876
rect 72940 56252 72996 56308
rect 71820 53340 71876 53396
rect 71148 53170 71204 53172
rect 71148 53118 71150 53170
rect 71150 53118 71202 53170
rect 71202 53118 71204 53170
rect 71148 53116 71204 53118
rect 72492 52892 72548 52948
rect 71260 52332 71316 52388
rect 71708 52220 71764 52276
rect 72828 52780 72884 52836
rect 72044 51436 72100 51492
rect 72268 51324 72324 51380
rect 68908 49922 68964 49924
rect 68908 49870 68910 49922
rect 68910 49870 68962 49922
rect 68962 49870 68964 49922
rect 68908 49868 68964 49870
rect 68796 48972 68852 49028
rect 67900 47964 67956 48020
rect 68348 47292 68404 47348
rect 67228 44156 67284 44212
rect 67228 42812 67284 42868
rect 67452 45052 67508 45108
rect 65436 41468 65492 41524
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65548 41298 65604 41300
rect 65548 41246 65550 41298
rect 65550 41246 65602 41298
rect 65602 41246 65604 41298
rect 65548 41244 65604 41246
rect 64540 37996 64596 38052
rect 64428 37324 64484 37380
rect 63756 35980 63812 36036
rect 64316 35980 64372 36036
rect 63308 34300 63364 34356
rect 63644 34972 63700 35028
rect 64988 37324 65044 37380
rect 65548 41020 65604 41076
rect 65996 41186 66052 41188
rect 65996 41134 65998 41186
rect 65998 41134 66050 41186
rect 66050 41134 66052 41186
rect 65996 41132 66052 41134
rect 66444 41132 66500 41188
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65660 38668 65716 38724
rect 68684 47852 68740 47908
rect 69692 49810 69748 49812
rect 69692 49758 69694 49810
rect 69694 49758 69746 49810
rect 69746 49758 69748 49810
rect 69692 49756 69748 49758
rect 69580 49026 69636 49028
rect 69580 48974 69582 49026
rect 69582 48974 69634 49026
rect 69634 48974 69636 49026
rect 69580 48972 69636 48974
rect 69356 47964 69412 48020
rect 68572 47346 68628 47348
rect 68572 47294 68574 47346
rect 68574 47294 68626 47346
rect 68626 47294 68628 47346
rect 68572 47292 68628 47294
rect 69580 47458 69636 47460
rect 69580 47406 69582 47458
rect 69582 47406 69634 47458
rect 69634 47406 69636 47458
rect 69580 47404 69636 47406
rect 68460 47068 68516 47124
rect 69244 47068 69300 47124
rect 69692 46562 69748 46564
rect 69692 46510 69694 46562
rect 69694 46510 69746 46562
rect 69746 46510 69748 46562
rect 69692 46508 69748 46510
rect 70700 50540 70756 50596
rect 71148 50594 71204 50596
rect 71148 50542 71150 50594
rect 71150 50542 71202 50594
rect 71202 50542 71204 50594
rect 71148 50540 71204 50542
rect 70028 49980 70084 50036
rect 69916 49196 69972 49252
rect 70476 50370 70532 50372
rect 70476 50318 70478 50370
rect 70478 50318 70530 50370
rect 70530 50318 70532 50370
rect 70476 50316 70532 50318
rect 70364 49810 70420 49812
rect 70364 49758 70366 49810
rect 70366 49758 70418 49810
rect 70418 49758 70420 49810
rect 70364 49756 70420 49758
rect 71708 50316 71764 50372
rect 72156 50034 72212 50036
rect 72156 49982 72158 50034
rect 72158 49982 72210 50034
rect 72210 49982 72212 50034
rect 72156 49980 72212 49982
rect 70588 49420 70644 49476
rect 70812 49420 70868 49476
rect 70028 47346 70084 47348
rect 70028 47294 70030 47346
rect 70030 47294 70082 47346
rect 70082 47294 70084 47346
rect 70028 47292 70084 47294
rect 70140 46562 70196 46564
rect 70140 46510 70142 46562
rect 70142 46510 70194 46562
rect 70194 46510 70196 46562
rect 70140 46508 70196 46510
rect 69468 45052 69524 45108
rect 68012 43820 68068 43876
rect 67676 41186 67732 41188
rect 67676 41134 67678 41186
rect 67678 41134 67730 41186
rect 67730 41134 67732 41186
rect 67676 41132 67732 41134
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65324 37996 65380 38052
rect 66556 37938 66612 37940
rect 66556 37886 66558 37938
rect 66558 37886 66610 37938
rect 66610 37886 66612 37938
rect 66556 37884 66612 37886
rect 67564 38050 67620 38052
rect 67564 37998 67566 38050
rect 67566 37998 67618 38050
rect 67618 37998 67620 38050
rect 67564 37996 67620 37998
rect 67228 37938 67284 37940
rect 67228 37886 67230 37938
rect 67230 37886 67282 37938
rect 67282 37886 67284 37938
rect 67228 37884 67284 37886
rect 65212 37324 65268 37380
rect 66780 37266 66836 37268
rect 66780 37214 66782 37266
rect 66782 37214 66834 37266
rect 66834 37214 66836 37266
rect 66780 37212 66836 37214
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 66108 34972 66164 35028
rect 63868 34860 63924 34916
rect 65324 34914 65380 34916
rect 65324 34862 65326 34914
rect 65326 34862 65378 34914
rect 65378 34862 65380 34914
rect 65324 34860 65380 34862
rect 64540 34354 64596 34356
rect 64540 34302 64542 34354
rect 64542 34302 64594 34354
rect 64594 34302 64596 34354
rect 64540 34300 64596 34302
rect 65884 34300 65940 34356
rect 69356 43426 69412 43428
rect 69356 43374 69358 43426
rect 69358 43374 69410 43426
rect 69410 43374 69412 43426
rect 69356 43372 69412 43374
rect 68572 42866 68628 42868
rect 68572 42814 68574 42866
rect 68574 42814 68626 42866
rect 68626 42814 68628 42866
rect 68572 42812 68628 42814
rect 69356 42812 69412 42868
rect 68684 41804 68740 41860
rect 69244 41858 69300 41860
rect 69244 41806 69246 41858
rect 69246 41806 69298 41858
rect 69298 41806 69300 41858
rect 69244 41804 69300 41806
rect 70364 47180 70420 47236
rect 70140 45052 70196 45108
rect 70028 43538 70084 43540
rect 70028 43486 70030 43538
rect 70030 43486 70082 43538
rect 70082 43486 70084 43538
rect 70028 43484 70084 43486
rect 70364 43372 70420 43428
rect 71484 49308 71540 49364
rect 71932 49308 71988 49364
rect 70812 47404 70868 47460
rect 71260 48636 71316 48692
rect 71596 48300 71652 48356
rect 71260 47234 71316 47236
rect 71260 47182 71262 47234
rect 71262 47182 71314 47234
rect 71314 47182 71316 47234
rect 71260 47180 71316 47182
rect 72492 50092 72548 50148
rect 72380 48412 72436 48468
rect 72268 48354 72324 48356
rect 72268 48302 72270 48354
rect 72270 48302 72322 48354
rect 72322 48302 72324 48354
rect 72268 48300 72324 48302
rect 70588 46898 70644 46900
rect 70588 46846 70590 46898
rect 70590 46846 70642 46898
rect 70642 46846 70644 46898
rect 70588 46844 70644 46846
rect 72268 47346 72324 47348
rect 72268 47294 72270 47346
rect 72270 47294 72322 47346
rect 72322 47294 72324 47346
rect 72268 47292 72324 47294
rect 72492 46732 72548 46788
rect 71260 44380 71316 44436
rect 70924 43538 70980 43540
rect 70924 43486 70926 43538
rect 70926 43486 70978 43538
rect 70978 43486 70980 43538
rect 70924 43484 70980 43486
rect 71484 43372 71540 43428
rect 72268 45052 72324 45108
rect 72268 44044 72324 44100
rect 72044 43650 72100 43652
rect 72044 43598 72046 43650
rect 72046 43598 72098 43650
rect 72098 43598 72100 43650
rect 72044 43596 72100 43598
rect 70476 41804 70532 41860
rect 70812 41804 70868 41860
rect 69468 41298 69524 41300
rect 69468 41246 69470 41298
rect 69470 41246 69522 41298
rect 69522 41246 69524 41298
rect 69468 41244 69524 41246
rect 68572 39004 68628 39060
rect 68236 38668 68292 38724
rect 68348 38108 68404 38164
rect 69692 39058 69748 39060
rect 69692 39006 69694 39058
rect 69694 39006 69746 39058
rect 69746 39006 69748 39058
rect 69692 39004 69748 39006
rect 69916 41132 69972 41188
rect 69916 40962 69972 40964
rect 69916 40910 69918 40962
rect 69918 40910 69970 40962
rect 69970 40910 69972 40962
rect 69916 40908 69972 40910
rect 70700 41580 70756 41636
rect 70364 41298 70420 41300
rect 70364 41246 70366 41298
rect 70366 41246 70418 41298
rect 70418 41246 70420 41298
rect 70364 41244 70420 41246
rect 71708 41916 71764 41972
rect 72380 44434 72436 44436
rect 72380 44382 72382 44434
rect 72382 44382 72434 44434
rect 72434 44382 72436 44434
rect 72380 44380 72436 44382
rect 72380 43708 72436 43764
rect 70924 41244 70980 41300
rect 70812 40908 70868 40964
rect 71260 41132 71316 41188
rect 71820 41186 71876 41188
rect 71820 41134 71822 41186
rect 71822 41134 71874 41186
rect 71874 41134 71876 41186
rect 71820 41132 71876 41134
rect 70252 39676 70308 39732
rect 70700 39730 70756 39732
rect 70700 39678 70702 39730
rect 70702 39678 70754 39730
rect 70754 39678 70756 39730
rect 70700 39676 70756 39678
rect 71260 39676 71316 39732
rect 70700 39004 70756 39060
rect 71372 39058 71428 39060
rect 71372 39006 71374 39058
rect 71374 39006 71426 39058
rect 71426 39006 71428 39058
rect 71372 39004 71428 39006
rect 69804 38668 69860 38724
rect 69244 38162 69300 38164
rect 69244 38110 69246 38162
rect 69246 38110 69298 38162
rect 69298 38110 69300 38162
rect 69244 38108 69300 38110
rect 68348 37660 68404 37716
rect 69580 37996 69636 38052
rect 66668 35586 66724 35588
rect 66668 35534 66670 35586
rect 66670 35534 66722 35586
rect 66722 35534 66724 35586
rect 66668 35532 66724 35534
rect 67228 35532 67284 35588
rect 66668 35026 66724 35028
rect 66668 34974 66670 35026
rect 66670 34974 66722 35026
rect 66722 34974 66724 35026
rect 66668 34972 66724 34974
rect 64988 34188 65044 34244
rect 63868 34018 63924 34020
rect 63868 33966 63870 34018
rect 63870 33966 63922 34018
rect 63922 33966 63924 34018
rect 63868 33964 63924 33966
rect 65772 34242 65828 34244
rect 65772 34190 65774 34242
rect 65774 34190 65826 34242
rect 65826 34190 65828 34242
rect 65772 34188 65828 34190
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 64988 33346 65044 33348
rect 64988 33294 64990 33346
rect 64990 33294 65042 33346
rect 65042 33294 65044 33346
rect 64988 33292 65044 33294
rect 65772 33346 65828 33348
rect 65772 33294 65774 33346
rect 65774 33294 65826 33346
rect 65826 33294 65828 33346
rect 65772 33292 65828 33294
rect 62636 32674 62692 32676
rect 62636 32622 62638 32674
rect 62638 32622 62690 32674
rect 62690 32622 62692 32674
rect 62636 32620 62692 32622
rect 66332 33292 66388 33348
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 66444 31612 66500 31668
rect 70140 37212 70196 37268
rect 68348 36370 68404 36372
rect 68348 36318 68350 36370
rect 68350 36318 68402 36370
rect 68402 36318 68404 36370
rect 68348 36316 68404 36318
rect 69468 36370 69524 36372
rect 69468 36318 69470 36370
rect 69470 36318 69522 36370
rect 69522 36318 69524 36370
rect 69468 36316 69524 36318
rect 68236 34860 68292 34916
rect 68460 34636 68516 34692
rect 68572 34860 68628 34916
rect 69692 34914 69748 34916
rect 69692 34862 69694 34914
rect 69694 34862 69746 34914
rect 69746 34862 69748 34914
rect 69692 34860 69748 34862
rect 69356 34690 69412 34692
rect 69356 34638 69358 34690
rect 69358 34638 69410 34690
rect 69410 34638 69412 34690
rect 69356 34636 69412 34638
rect 70588 36764 70644 36820
rect 70364 36370 70420 36372
rect 70364 36318 70366 36370
rect 70366 36318 70418 36370
rect 70418 36318 70420 36370
rect 70364 36316 70420 36318
rect 68684 33292 68740 33348
rect 67676 32396 67732 32452
rect 68572 32450 68628 32452
rect 68572 32398 68574 32450
rect 68574 32398 68626 32450
rect 68626 32398 68628 32450
rect 68572 32396 68628 32398
rect 67452 31724 67508 31780
rect 68012 32284 68068 32340
rect 69692 33346 69748 33348
rect 69692 33294 69694 33346
rect 69694 33294 69746 33346
rect 69746 33294 69748 33346
rect 69692 33292 69748 33294
rect 71148 36764 71204 36820
rect 72268 41580 72324 41636
rect 72268 41356 72324 41412
rect 72268 41020 72324 41076
rect 72044 40348 72100 40404
rect 71932 39004 71988 39060
rect 71708 36764 71764 36820
rect 70812 36316 70868 36372
rect 72716 48412 72772 48468
rect 72828 47292 72884 47348
rect 74956 66162 75012 66164
rect 74956 66110 74958 66162
rect 74958 66110 75010 66162
rect 75010 66110 75012 66162
rect 74956 66108 75012 66110
rect 74956 64652 75012 64708
rect 74956 63868 75012 63924
rect 74396 62748 74452 62804
rect 74732 62748 74788 62804
rect 74508 62412 74564 62468
rect 74396 61964 74452 62020
rect 74284 61852 74340 61908
rect 74508 60002 74564 60004
rect 74508 59950 74510 60002
rect 74510 59950 74562 60002
rect 74562 59950 74564 60002
rect 74508 59948 74564 59950
rect 73724 59500 73780 59556
rect 73500 59276 73556 59332
rect 73612 58380 73668 58436
rect 74172 58380 74228 58436
rect 74284 58492 74340 58548
rect 74060 58268 74116 58324
rect 73388 57596 73444 57652
rect 74060 58044 74116 58100
rect 74172 57820 74228 57876
rect 73724 57596 73780 57652
rect 74060 56924 74116 56980
rect 73500 56194 73556 56196
rect 73500 56142 73502 56194
rect 73502 56142 73554 56194
rect 73554 56142 73556 56194
rect 73500 56140 73556 56142
rect 74620 58940 74676 58996
rect 74620 58268 74676 58324
rect 74844 62466 74900 62468
rect 74844 62414 74846 62466
rect 74846 62414 74898 62466
rect 74898 62414 74900 62466
rect 74844 62412 74900 62414
rect 75292 67676 75348 67732
rect 75516 67900 75572 67956
rect 75404 67618 75460 67620
rect 75404 67566 75406 67618
rect 75406 67566 75458 67618
rect 75458 67566 75460 67618
rect 75404 67564 75460 67566
rect 75516 67228 75572 67284
rect 76300 68626 76356 68628
rect 76300 68574 76302 68626
rect 76302 68574 76354 68626
rect 76354 68574 76356 68626
rect 76300 68572 76356 68574
rect 75740 67116 75796 67172
rect 75516 66892 75572 66948
rect 75964 66332 76020 66388
rect 75404 65324 75460 65380
rect 75404 63868 75460 63924
rect 75740 65884 75796 65940
rect 75180 63644 75236 63700
rect 75740 63644 75796 63700
rect 75404 63532 75460 63588
rect 75516 63420 75572 63476
rect 75404 62354 75460 62356
rect 75404 62302 75406 62354
rect 75406 62302 75458 62354
rect 75458 62302 75460 62354
rect 75404 62300 75460 62302
rect 75404 62076 75460 62132
rect 75404 61628 75460 61684
rect 75180 61292 75236 61348
rect 74284 57650 74340 57652
rect 74284 57598 74286 57650
rect 74286 57598 74338 57650
rect 74338 57598 74340 57650
rect 74284 57596 74340 57598
rect 74844 59388 74900 59444
rect 74172 56588 74228 56644
rect 75068 57708 75124 57764
rect 74956 57148 75012 57204
rect 74732 57036 74788 57092
rect 73948 56306 74004 56308
rect 73948 56254 73950 56306
rect 73950 56254 74002 56306
rect 74002 56254 74004 56306
rect 73948 56252 74004 56254
rect 74844 56924 74900 56980
rect 73836 56140 73892 56196
rect 73388 55356 73444 55412
rect 74060 54684 74116 54740
rect 73500 53564 73556 53620
rect 73500 52274 73556 52276
rect 73500 52222 73502 52274
rect 73502 52222 73554 52274
rect 73554 52222 73556 52274
rect 73500 52220 73556 52222
rect 73836 52892 73892 52948
rect 73948 52332 74004 52388
rect 73724 51884 73780 51940
rect 74060 51996 74116 52052
rect 73276 51378 73332 51380
rect 73276 51326 73278 51378
rect 73278 51326 73330 51378
rect 73330 51326 73332 51378
rect 73276 51324 73332 51326
rect 73500 51490 73556 51492
rect 73500 51438 73502 51490
rect 73502 51438 73554 51490
rect 73554 51438 73556 51490
rect 73500 51436 73556 51438
rect 73948 51436 74004 51492
rect 73612 51378 73668 51380
rect 73612 51326 73614 51378
rect 73614 51326 73666 51378
rect 73666 51326 73668 51378
rect 73612 51324 73668 51326
rect 73388 50092 73444 50148
rect 73612 51100 73668 51156
rect 73612 50540 73668 50596
rect 73388 49922 73444 49924
rect 73388 49870 73390 49922
rect 73390 49870 73442 49922
rect 73442 49870 73444 49922
rect 73388 49868 73444 49870
rect 73052 47628 73108 47684
rect 73724 50428 73780 50484
rect 73836 48130 73892 48132
rect 73836 48078 73838 48130
rect 73838 48078 73890 48130
rect 73890 48078 73892 48130
rect 73836 48076 73892 48078
rect 72828 44098 72884 44100
rect 72828 44046 72830 44098
rect 72830 44046 72882 44098
rect 72882 44046 72884 44098
rect 72828 44044 72884 44046
rect 72716 43650 72772 43652
rect 72716 43598 72718 43650
rect 72718 43598 72770 43650
rect 72770 43598 72772 43650
rect 72716 43596 72772 43598
rect 73612 47628 73668 47684
rect 73388 47292 73444 47348
rect 73164 46844 73220 46900
rect 73164 45948 73220 46004
rect 73276 42476 73332 42532
rect 73276 41970 73332 41972
rect 73276 41918 73278 41970
rect 73278 41918 73330 41970
rect 73330 41918 73332 41970
rect 73276 41916 73332 41918
rect 73948 46898 74004 46900
rect 73948 46846 73950 46898
rect 73950 46846 74002 46898
rect 74002 46846 74004 46898
rect 73948 46844 74004 46846
rect 73836 46786 73892 46788
rect 73836 46734 73838 46786
rect 73838 46734 73890 46786
rect 73890 46734 73892 46786
rect 73836 46732 73892 46734
rect 74956 56364 75012 56420
rect 74956 55468 75012 55524
rect 74844 55356 74900 55412
rect 74956 54738 75012 54740
rect 74956 54686 74958 54738
rect 74958 54686 75010 54738
rect 75010 54686 75012 54738
rect 74956 54684 75012 54686
rect 74396 53676 74452 53732
rect 74396 52834 74452 52836
rect 74396 52782 74398 52834
rect 74398 52782 74450 52834
rect 74450 52782 74452 52834
rect 74396 52780 74452 52782
rect 74508 51602 74564 51604
rect 74508 51550 74510 51602
rect 74510 51550 74562 51602
rect 74562 51550 74564 51602
rect 74508 51548 74564 51550
rect 74284 50316 74340 50372
rect 74844 53900 74900 53956
rect 74732 53116 74788 53172
rect 74732 51996 74788 52052
rect 75292 60396 75348 60452
rect 76188 65884 76244 65940
rect 76076 65548 76132 65604
rect 75964 63756 76020 63812
rect 75964 63196 76020 63252
rect 76076 63308 76132 63364
rect 75852 62636 75908 62692
rect 75628 62300 75684 62356
rect 75740 62076 75796 62132
rect 75628 61570 75684 61572
rect 75628 61518 75630 61570
rect 75630 61518 75682 61570
rect 75682 61518 75684 61570
rect 75628 61516 75684 61518
rect 75292 57932 75348 57988
rect 76412 63868 76468 63924
rect 78540 73500 78596 73556
rect 76636 71650 76692 71652
rect 76636 71598 76638 71650
rect 76638 71598 76690 71650
rect 76690 71598 76692 71650
rect 76636 71596 76692 71598
rect 76972 69132 77028 69188
rect 77196 70028 77252 70084
rect 77420 69298 77476 69300
rect 77420 69246 77422 69298
rect 77422 69246 77474 69298
rect 77474 69246 77476 69298
rect 77420 69244 77476 69246
rect 78316 70082 78372 70084
rect 78316 70030 78318 70082
rect 78318 70030 78370 70082
rect 78370 70030 78372 70082
rect 78316 70028 78372 70030
rect 78876 77420 78932 77476
rect 78764 76972 78820 77028
rect 78764 76076 78820 76132
rect 79884 78988 79940 79044
rect 79436 77308 79492 77364
rect 79212 77196 79268 77252
rect 79212 76972 79268 77028
rect 80332 81900 80388 81956
rect 80444 82236 80500 82292
rect 80668 82236 80724 82292
rect 81276 83130 81332 83132
rect 81276 83078 81278 83130
rect 81278 83078 81330 83130
rect 81330 83078 81332 83130
rect 81276 83076 81332 83078
rect 81380 83130 81436 83132
rect 81380 83078 81382 83130
rect 81382 83078 81434 83130
rect 81434 83078 81436 83130
rect 81380 83076 81436 83078
rect 81484 83130 81540 83132
rect 81484 83078 81486 83130
rect 81486 83078 81538 83130
rect 81538 83078 81540 83130
rect 81484 83076 81540 83078
rect 81452 82236 81508 82292
rect 96636 94890 96692 94892
rect 96636 94838 96638 94890
rect 96638 94838 96690 94890
rect 96690 94838 96692 94890
rect 96636 94836 96692 94838
rect 96740 94890 96796 94892
rect 96740 94838 96742 94890
rect 96742 94838 96794 94890
rect 96794 94838 96796 94890
rect 96740 94836 96796 94838
rect 96844 94890 96900 94892
rect 96844 94838 96846 94890
rect 96846 94838 96898 94890
rect 96898 94838 96900 94890
rect 96844 94836 96900 94838
rect 96636 93322 96692 93324
rect 96636 93270 96638 93322
rect 96638 93270 96690 93322
rect 96690 93270 96692 93322
rect 96636 93268 96692 93270
rect 96740 93322 96796 93324
rect 96740 93270 96742 93322
rect 96742 93270 96794 93322
rect 96794 93270 96796 93322
rect 96740 93268 96796 93270
rect 96844 93322 96900 93324
rect 96844 93270 96846 93322
rect 96846 93270 96898 93322
rect 96898 93270 96900 93322
rect 96844 93268 96900 93270
rect 96636 91754 96692 91756
rect 96636 91702 96638 91754
rect 96638 91702 96690 91754
rect 96690 91702 96692 91754
rect 96636 91700 96692 91702
rect 96740 91754 96796 91756
rect 96740 91702 96742 91754
rect 96742 91702 96794 91754
rect 96794 91702 96796 91754
rect 96740 91700 96796 91702
rect 96844 91754 96900 91756
rect 96844 91702 96846 91754
rect 96846 91702 96898 91754
rect 96898 91702 96900 91754
rect 96844 91700 96900 91702
rect 96636 90186 96692 90188
rect 96636 90134 96638 90186
rect 96638 90134 96690 90186
rect 96690 90134 96692 90186
rect 96636 90132 96692 90134
rect 96740 90186 96796 90188
rect 96740 90134 96742 90186
rect 96742 90134 96794 90186
rect 96794 90134 96796 90186
rect 96740 90132 96796 90134
rect 96844 90186 96900 90188
rect 96844 90134 96846 90186
rect 96846 90134 96898 90186
rect 96898 90134 96900 90186
rect 96844 90132 96900 90134
rect 87052 86828 87108 86884
rect 82348 85708 82404 85764
rect 85596 86492 85652 86548
rect 82460 86380 82516 86436
rect 82124 84194 82180 84196
rect 82124 84142 82126 84194
rect 82126 84142 82178 84194
rect 82178 84142 82180 84194
rect 82124 84140 82180 84142
rect 82012 83356 82068 83412
rect 82012 82572 82068 82628
rect 80444 81340 80500 81396
rect 80556 81452 80612 81508
rect 80444 81116 80500 81172
rect 80332 80780 80388 80836
rect 80668 81228 80724 81284
rect 80556 81004 80612 81060
rect 81276 81562 81332 81564
rect 81276 81510 81278 81562
rect 81278 81510 81330 81562
rect 81330 81510 81332 81562
rect 81276 81508 81332 81510
rect 81380 81562 81436 81564
rect 81380 81510 81382 81562
rect 81382 81510 81434 81562
rect 81434 81510 81436 81562
rect 81380 81508 81436 81510
rect 81484 81562 81540 81564
rect 81484 81510 81486 81562
rect 81486 81510 81538 81562
rect 81538 81510 81540 81562
rect 81484 81508 81540 81510
rect 81116 80556 81172 80612
rect 81676 81228 81732 81284
rect 81564 81170 81620 81172
rect 81564 81118 81566 81170
rect 81566 81118 81618 81170
rect 81618 81118 81620 81170
rect 81564 81116 81620 81118
rect 81452 80946 81508 80948
rect 81452 80894 81454 80946
rect 81454 80894 81506 80946
rect 81506 80894 81508 80946
rect 81452 80892 81508 80894
rect 81340 80220 81396 80276
rect 81276 79994 81332 79996
rect 81276 79942 81278 79994
rect 81278 79942 81330 79994
rect 81330 79942 81332 79994
rect 81276 79940 81332 79942
rect 81380 79994 81436 79996
rect 81380 79942 81382 79994
rect 81382 79942 81434 79994
rect 81434 79942 81436 79994
rect 81380 79940 81436 79942
rect 81484 79994 81540 79996
rect 81484 79942 81486 79994
rect 81486 79942 81538 79994
rect 81538 79942 81540 79994
rect 81484 79940 81540 79942
rect 80668 79714 80724 79716
rect 80668 79662 80670 79714
rect 80670 79662 80722 79714
rect 80722 79662 80724 79714
rect 80668 79660 80724 79662
rect 81452 79602 81508 79604
rect 81452 79550 81454 79602
rect 81454 79550 81506 79602
rect 81506 79550 81508 79602
rect 81452 79548 81508 79550
rect 80444 78988 80500 79044
rect 82348 81282 82404 81284
rect 82348 81230 82350 81282
rect 82350 81230 82402 81282
rect 82402 81230 82404 81282
rect 82348 81228 82404 81230
rect 82124 81170 82180 81172
rect 82124 81118 82126 81170
rect 82126 81118 82178 81170
rect 82178 81118 82180 81170
rect 82124 81116 82180 81118
rect 82572 85090 82628 85092
rect 82572 85038 82574 85090
rect 82574 85038 82626 85090
rect 82626 85038 82628 85090
rect 82572 85036 82628 85038
rect 83132 86434 83188 86436
rect 83132 86382 83134 86434
rect 83134 86382 83186 86434
rect 83186 86382 83188 86434
rect 83132 86380 83188 86382
rect 82796 85596 82852 85652
rect 83468 85036 83524 85092
rect 82684 84028 82740 84084
rect 83020 84252 83076 84308
rect 83020 82236 83076 82292
rect 82684 81954 82740 81956
rect 82684 81902 82686 81954
rect 82686 81902 82738 81954
rect 82738 81902 82740 81954
rect 82684 81900 82740 81902
rect 87052 86434 87108 86436
rect 87052 86382 87054 86434
rect 87054 86382 87106 86434
rect 87106 86382 87108 86434
rect 87052 86380 87108 86382
rect 88396 87500 88452 87556
rect 87612 86882 87668 86884
rect 87612 86830 87614 86882
rect 87614 86830 87666 86882
rect 87666 86830 87668 86882
rect 87612 86828 87668 86830
rect 88172 86380 88228 86436
rect 87948 86268 88004 86324
rect 87276 85932 87332 85988
rect 87724 85986 87780 85988
rect 87724 85934 87726 85986
rect 87726 85934 87778 85986
rect 87778 85934 87780 85986
rect 87724 85932 87780 85934
rect 89516 87554 89572 87556
rect 89516 87502 89518 87554
rect 89518 87502 89570 87554
rect 89570 87502 89572 87554
rect 89516 87500 89572 87502
rect 90860 87500 90916 87556
rect 88732 86546 88788 86548
rect 88732 86494 88734 86546
rect 88734 86494 88786 86546
rect 88786 86494 88788 86546
rect 88732 86492 88788 86494
rect 89740 86492 89796 86548
rect 89180 86380 89236 86436
rect 86492 85260 86548 85316
rect 88060 85708 88116 85764
rect 87500 85148 87556 85204
rect 84924 84418 84980 84420
rect 84924 84366 84926 84418
rect 84926 84366 84978 84418
rect 84978 84366 84980 84418
rect 84924 84364 84980 84366
rect 83580 83410 83636 83412
rect 83580 83358 83582 83410
rect 83582 83358 83634 83410
rect 83634 83358 83636 83410
rect 83580 83356 83636 83358
rect 83468 82236 83524 82292
rect 82908 81564 82964 81620
rect 82460 81004 82516 81060
rect 82908 80780 82964 80836
rect 81788 78988 81844 79044
rect 81276 78426 81332 78428
rect 81276 78374 81278 78426
rect 81278 78374 81330 78426
rect 81330 78374 81332 78426
rect 81276 78372 81332 78374
rect 81380 78426 81436 78428
rect 81380 78374 81382 78426
rect 81382 78374 81434 78426
rect 81434 78374 81436 78426
rect 81380 78372 81436 78374
rect 81484 78426 81540 78428
rect 81484 78374 81486 78426
rect 81486 78374 81538 78426
rect 81538 78374 81540 78426
rect 81484 78372 81540 78374
rect 81340 77868 81396 77924
rect 80780 77308 80836 77364
rect 80444 77250 80500 77252
rect 80444 77198 80446 77250
rect 80446 77198 80498 77250
rect 80498 77198 80500 77250
rect 80444 77196 80500 77198
rect 82012 80668 82068 80724
rect 82908 80386 82964 80388
rect 82908 80334 82910 80386
rect 82910 80334 82962 80386
rect 82962 80334 82964 80386
rect 82908 80332 82964 80334
rect 83020 80220 83076 80276
rect 82236 80162 82292 80164
rect 82236 80110 82238 80162
rect 82238 80110 82290 80162
rect 82290 80110 82292 80162
rect 82236 80108 82292 80110
rect 82124 79714 82180 79716
rect 82124 79662 82126 79714
rect 82126 79662 82178 79714
rect 82178 79662 82180 79714
rect 82124 79660 82180 79662
rect 82124 77922 82180 77924
rect 82124 77870 82126 77922
rect 82126 77870 82178 77922
rect 82178 77870 82180 77922
rect 82124 77868 82180 77870
rect 82796 78764 82852 78820
rect 83692 81730 83748 81732
rect 83692 81678 83694 81730
rect 83694 81678 83746 81730
rect 83746 81678 83748 81730
rect 83692 81676 83748 81678
rect 83692 81058 83748 81060
rect 83692 81006 83694 81058
rect 83694 81006 83746 81058
rect 83746 81006 83748 81058
rect 83692 81004 83748 81006
rect 83580 80610 83636 80612
rect 83580 80558 83582 80610
rect 83582 80558 83634 80610
rect 83634 80558 83636 80610
rect 83580 80556 83636 80558
rect 83580 80274 83636 80276
rect 83580 80222 83582 80274
rect 83582 80222 83634 80274
rect 83634 80222 83636 80274
rect 83580 80220 83636 80222
rect 83132 79436 83188 79492
rect 83244 80108 83300 80164
rect 83132 79212 83188 79268
rect 83020 77138 83076 77140
rect 83020 77086 83022 77138
rect 83022 77086 83074 77138
rect 83074 77086 83076 77138
rect 83020 77084 83076 77086
rect 81276 76858 81332 76860
rect 81276 76806 81278 76858
rect 81278 76806 81330 76858
rect 81330 76806 81332 76858
rect 81276 76804 81332 76806
rect 81380 76858 81436 76860
rect 81380 76806 81382 76858
rect 81382 76806 81434 76858
rect 81434 76806 81436 76858
rect 81380 76804 81436 76806
rect 81484 76858 81540 76860
rect 81484 76806 81486 76858
rect 81486 76806 81538 76858
rect 81538 76806 81540 76858
rect 81484 76804 81540 76806
rect 80780 76636 80836 76692
rect 80556 76412 80612 76468
rect 79772 75794 79828 75796
rect 79772 75742 79774 75794
rect 79774 75742 79826 75794
rect 79826 75742 79828 75794
rect 79772 75740 79828 75742
rect 81228 75740 81284 75796
rect 81564 76188 81620 76244
rect 82796 76578 82852 76580
rect 82796 76526 82798 76578
rect 82798 76526 82850 76578
rect 82850 76526 82852 76578
rect 82796 76524 82852 76526
rect 82348 76466 82404 76468
rect 82348 76414 82350 76466
rect 82350 76414 82402 76466
rect 82402 76414 82404 76466
rect 82348 76412 82404 76414
rect 82236 76242 82292 76244
rect 82236 76190 82238 76242
rect 82238 76190 82290 76242
rect 82290 76190 82292 76242
rect 82236 76188 82292 76190
rect 81452 75628 81508 75684
rect 82348 75682 82404 75684
rect 82348 75630 82350 75682
rect 82350 75630 82402 75682
rect 82402 75630 82404 75682
rect 82348 75628 82404 75630
rect 83468 79212 83524 79268
rect 83580 79548 83636 79604
rect 83580 78876 83636 78932
rect 83356 78706 83412 78708
rect 83356 78654 83358 78706
rect 83358 78654 83410 78706
rect 83410 78654 83412 78706
rect 83356 78652 83412 78654
rect 83356 77026 83412 77028
rect 83356 76974 83358 77026
rect 83358 76974 83410 77026
rect 83410 76974 83412 77026
rect 83356 76972 83412 76974
rect 83916 82684 83972 82740
rect 84140 82236 84196 82292
rect 84924 84082 84980 84084
rect 84924 84030 84926 84082
rect 84926 84030 84978 84082
rect 84978 84030 84980 84082
rect 84924 84028 84980 84030
rect 84252 81564 84308 81620
rect 84364 81004 84420 81060
rect 84140 80668 84196 80724
rect 84252 80386 84308 80388
rect 84252 80334 84254 80386
rect 84254 80334 84306 80386
rect 84306 80334 84308 80386
rect 84252 80332 84308 80334
rect 85036 82684 85092 82740
rect 84812 81676 84868 81732
rect 84588 81058 84644 81060
rect 84588 81006 84590 81058
rect 84590 81006 84642 81058
rect 84642 81006 84644 81058
rect 84588 81004 84644 81006
rect 85596 83692 85652 83748
rect 87388 83692 87444 83748
rect 85260 82626 85316 82628
rect 85260 82574 85262 82626
rect 85262 82574 85314 82626
rect 85314 82574 85316 82626
rect 85260 82572 85316 82574
rect 85260 81564 85316 81620
rect 86604 82626 86660 82628
rect 86604 82574 86606 82626
rect 86606 82574 86658 82626
rect 86658 82574 86660 82626
rect 86604 82572 86660 82574
rect 84476 80220 84532 80276
rect 84700 80220 84756 80276
rect 84364 79548 84420 79604
rect 84252 79490 84308 79492
rect 84252 79438 84254 79490
rect 84254 79438 84306 79490
rect 84306 79438 84308 79490
rect 84252 79436 84308 79438
rect 83692 78652 83748 78708
rect 84252 78764 84308 78820
rect 84140 78706 84196 78708
rect 84140 78654 84142 78706
rect 84142 78654 84194 78706
rect 84194 78654 84196 78706
rect 84140 78652 84196 78654
rect 85372 80332 85428 80388
rect 85260 79436 85316 79492
rect 84588 78092 84644 78148
rect 84364 77308 84420 77364
rect 85260 77196 85316 77252
rect 84700 77084 84756 77140
rect 82796 75628 82852 75684
rect 80556 75516 80612 75572
rect 82236 75404 82292 75460
rect 81276 75290 81332 75292
rect 81276 75238 81278 75290
rect 81278 75238 81330 75290
rect 81330 75238 81332 75290
rect 81276 75236 81332 75238
rect 81380 75290 81436 75292
rect 81380 75238 81382 75290
rect 81382 75238 81434 75290
rect 81434 75238 81436 75290
rect 81380 75236 81436 75238
rect 81484 75290 81540 75292
rect 81484 75238 81486 75290
rect 81486 75238 81538 75290
rect 81538 75238 81540 75290
rect 81484 75236 81540 75238
rect 78764 73442 78820 73444
rect 78764 73390 78766 73442
rect 78766 73390 78818 73442
rect 78818 73390 78820 73442
rect 78764 73388 78820 73390
rect 78652 69692 78708 69748
rect 77420 67676 77476 67732
rect 77084 67004 77140 67060
rect 76748 66892 76804 66948
rect 77420 66444 77476 66500
rect 76524 63420 76580 63476
rect 76860 64428 76916 64484
rect 76300 61852 76356 61908
rect 75852 60114 75908 60116
rect 75852 60062 75854 60114
rect 75854 60062 75906 60114
rect 75906 60062 75908 60114
rect 75852 60060 75908 60062
rect 75852 59052 75908 59108
rect 75628 58434 75684 58436
rect 75628 58382 75630 58434
rect 75630 58382 75682 58434
rect 75682 58382 75684 58434
rect 75628 58380 75684 58382
rect 75516 58044 75572 58100
rect 75404 57708 75460 57764
rect 75852 57762 75908 57764
rect 75852 57710 75854 57762
rect 75854 57710 75906 57762
rect 75906 57710 75908 57762
rect 75852 57708 75908 57710
rect 75292 57036 75348 57092
rect 76300 61180 76356 61236
rect 76524 62860 76580 62916
rect 76860 62524 76916 62580
rect 77084 63980 77140 64036
rect 77196 63868 77252 63924
rect 77308 63250 77364 63252
rect 77308 63198 77310 63250
rect 77310 63198 77362 63250
rect 77362 63198 77364 63250
rect 77308 63196 77364 63198
rect 77308 61570 77364 61572
rect 77308 61518 77310 61570
rect 77310 61518 77362 61570
rect 77362 61518 77364 61570
rect 77308 61516 77364 61518
rect 76972 61404 77028 61460
rect 76748 60674 76804 60676
rect 76748 60622 76750 60674
rect 76750 60622 76802 60674
rect 76802 60622 76804 60674
rect 76748 60620 76804 60622
rect 77644 66220 77700 66276
rect 78204 69244 78260 69300
rect 78540 69186 78596 69188
rect 78540 69134 78542 69186
rect 78542 69134 78594 69186
rect 78594 69134 78596 69186
rect 78540 69132 78596 69134
rect 78988 73106 79044 73108
rect 78988 73054 78990 73106
rect 78990 73054 79042 73106
rect 79042 73054 79044 73106
rect 78988 73052 79044 73054
rect 78988 72156 79044 72212
rect 79100 72268 79156 72324
rect 79100 69410 79156 69412
rect 79100 69358 79102 69410
rect 79102 69358 79154 69410
rect 79154 69358 79156 69410
rect 79100 69356 79156 69358
rect 79324 73554 79380 73556
rect 79324 73502 79326 73554
rect 79326 73502 79378 73554
rect 79378 73502 79380 73554
rect 79324 73500 79380 73502
rect 79996 73052 80052 73108
rect 79996 71596 80052 71652
rect 80332 72156 80388 72212
rect 82572 75458 82628 75460
rect 82572 75406 82574 75458
rect 82574 75406 82626 75458
rect 82626 75406 82628 75458
rect 82572 75404 82628 75406
rect 82236 74226 82292 74228
rect 82236 74174 82238 74226
rect 82238 74174 82290 74226
rect 82290 74174 82292 74226
rect 82236 74172 82292 74174
rect 83244 75516 83300 75572
rect 83020 74508 83076 74564
rect 82796 74172 82852 74228
rect 81276 73722 81332 73724
rect 81276 73670 81278 73722
rect 81278 73670 81330 73722
rect 81330 73670 81332 73722
rect 81276 73668 81332 73670
rect 81380 73722 81436 73724
rect 81380 73670 81382 73722
rect 81382 73670 81434 73722
rect 81434 73670 81436 73722
rect 81380 73668 81436 73670
rect 81484 73722 81540 73724
rect 81484 73670 81486 73722
rect 81486 73670 81538 73722
rect 81538 73670 81540 73722
rect 81484 73668 81540 73670
rect 81116 72156 81172 72212
rect 81276 72154 81332 72156
rect 81276 72102 81278 72154
rect 81278 72102 81330 72154
rect 81330 72102 81332 72154
rect 81276 72100 81332 72102
rect 81380 72154 81436 72156
rect 81380 72102 81382 72154
rect 81382 72102 81434 72154
rect 81434 72102 81436 72154
rect 81380 72100 81436 72102
rect 81484 72154 81540 72156
rect 81484 72102 81486 72154
rect 81486 72102 81538 72154
rect 81538 72102 81540 72154
rect 81484 72100 81540 72102
rect 80556 71650 80612 71652
rect 80556 71598 80558 71650
rect 80558 71598 80610 71650
rect 80610 71598 80612 71650
rect 80556 71596 80612 71598
rect 81564 71596 81620 71652
rect 82348 71202 82404 71204
rect 82348 71150 82350 71202
rect 82350 71150 82402 71202
rect 82402 71150 82404 71202
rect 82348 71148 82404 71150
rect 83468 75682 83524 75684
rect 83468 75630 83470 75682
rect 83470 75630 83522 75682
rect 83522 75630 83524 75682
rect 83468 75628 83524 75630
rect 84252 77026 84308 77028
rect 84252 76974 84254 77026
rect 84254 76974 84306 77026
rect 84306 76974 84308 77026
rect 84252 76972 84308 76974
rect 85596 80332 85652 80388
rect 85596 79996 85652 80052
rect 85484 79548 85540 79604
rect 85820 79996 85876 80052
rect 85372 76860 85428 76916
rect 85596 77308 85652 77364
rect 84028 75404 84084 75460
rect 84252 76300 84308 76356
rect 85372 76300 85428 76356
rect 84252 75628 84308 75684
rect 83580 74508 83636 74564
rect 83020 71820 83076 71876
rect 81452 70754 81508 70756
rect 81452 70702 81454 70754
rect 81454 70702 81506 70754
rect 81506 70702 81508 70754
rect 81452 70700 81508 70702
rect 81276 70586 81332 70588
rect 81276 70534 81278 70586
rect 81278 70534 81330 70586
rect 81330 70534 81332 70586
rect 81276 70532 81332 70534
rect 81380 70586 81436 70588
rect 81380 70534 81382 70586
rect 81382 70534 81434 70586
rect 81434 70534 81436 70586
rect 81380 70532 81436 70534
rect 81484 70586 81540 70588
rect 81484 70534 81486 70586
rect 81486 70534 81538 70586
rect 81538 70534 81540 70586
rect 81484 70532 81540 70534
rect 79996 69244 80052 69300
rect 78092 68738 78148 68740
rect 78092 68686 78094 68738
rect 78094 68686 78146 68738
rect 78146 68686 78148 68738
rect 78092 68684 78148 68686
rect 77980 68572 78036 68628
rect 77980 68012 78036 68068
rect 77756 66108 77812 66164
rect 77532 65884 77588 65940
rect 77868 65996 77924 66052
rect 78652 66332 78708 66388
rect 78540 66274 78596 66276
rect 78540 66222 78542 66274
rect 78542 66222 78594 66274
rect 78594 66222 78596 66274
rect 78540 66220 78596 66222
rect 78092 64988 78148 65044
rect 77868 64482 77924 64484
rect 77868 64430 77870 64482
rect 77870 64430 77922 64482
rect 77922 64430 77924 64482
rect 77868 64428 77924 64430
rect 77756 64092 77812 64148
rect 78428 65436 78484 65492
rect 78540 65772 78596 65828
rect 78540 65324 78596 65380
rect 78316 64540 78372 64596
rect 77980 63922 78036 63924
rect 77980 63870 77982 63922
rect 77982 63870 78034 63922
rect 78034 63870 78036 63922
rect 77980 63868 78036 63870
rect 77756 63308 77812 63364
rect 77868 63644 77924 63700
rect 77420 61292 77476 61348
rect 81228 69522 81284 69524
rect 81228 69470 81230 69522
rect 81230 69470 81282 69522
rect 81282 69470 81284 69522
rect 81228 69468 81284 69470
rect 79100 68684 79156 68740
rect 79100 67564 79156 67620
rect 79212 66892 79268 66948
rect 79324 68348 79380 68404
rect 79100 66556 79156 66612
rect 79100 65714 79156 65716
rect 79100 65662 79102 65714
rect 79102 65662 79154 65714
rect 79154 65662 79156 65714
rect 79100 65660 79156 65662
rect 79996 68402 80052 68404
rect 79996 68350 79998 68402
rect 79998 68350 80050 68402
rect 80050 68350 80052 68402
rect 79996 68348 80052 68350
rect 80108 67116 80164 67172
rect 81276 69018 81332 69020
rect 81276 68966 81278 69018
rect 81278 68966 81330 69018
rect 81330 68966 81332 69018
rect 81276 68964 81332 68966
rect 81380 69018 81436 69020
rect 81380 68966 81382 69018
rect 81382 68966 81434 69018
rect 81434 68966 81436 69018
rect 81380 68964 81436 68966
rect 81484 69018 81540 69020
rect 81484 68966 81486 69018
rect 81486 68966 81538 69018
rect 81538 68966 81540 69018
rect 81484 68964 81540 68966
rect 81276 67450 81332 67452
rect 81276 67398 81278 67450
rect 81278 67398 81330 67450
rect 81330 67398 81332 67450
rect 81276 67396 81332 67398
rect 81380 67450 81436 67452
rect 81380 67398 81382 67450
rect 81382 67398 81434 67450
rect 81434 67398 81436 67450
rect 81380 67396 81436 67398
rect 81484 67450 81540 67452
rect 81484 67398 81486 67450
rect 81486 67398 81538 67450
rect 81538 67398 81540 67450
rect 81484 67396 81540 67398
rect 81228 67170 81284 67172
rect 81228 67118 81230 67170
rect 81230 67118 81282 67170
rect 81282 67118 81284 67170
rect 81228 67116 81284 67118
rect 80556 66946 80612 66948
rect 80556 66894 80558 66946
rect 80558 66894 80610 66946
rect 80610 66894 80612 66946
rect 80556 66892 80612 66894
rect 79660 65602 79716 65604
rect 79660 65550 79662 65602
rect 79662 65550 79714 65602
rect 79714 65550 79716 65602
rect 79660 65548 79716 65550
rect 80668 66780 80724 66836
rect 80668 65884 80724 65940
rect 79996 65490 80052 65492
rect 79996 65438 79998 65490
rect 79998 65438 80050 65490
rect 80050 65438 80052 65490
rect 79996 65436 80052 65438
rect 79660 65100 79716 65156
rect 78988 64876 79044 64932
rect 79436 64988 79492 65044
rect 78988 64594 79044 64596
rect 78988 64542 78990 64594
rect 78990 64542 79042 64594
rect 79042 64542 79044 64594
rect 78988 64540 79044 64542
rect 79100 64092 79156 64148
rect 79324 64316 79380 64372
rect 78764 63756 78820 63812
rect 78540 63138 78596 63140
rect 78540 63086 78542 63138
rect 78542 63086 78594 63138
rect 78594 63086 78596 63138
rect 78540 63084 78596 63086
rect 77980 61404 78036 61460
rect 78764 63026 78820 63028
rect 78764 62974 78766 63026
rect 78766 62974 78818 63026
rect 78818 62974 78820 63026
rect 78764 62972 78820 62974
rect 78092 62076 78148 62132
rect 77868 60956 77924 61012
rect 77532 60396 77588 60452
rect 76972 60172 77028 60228
rect 77644 60172 77700 60228
rect 76524 60060 76580 60116
rect 76188 58940 76244 58996
rect 76076 58492 76132 58548
rect 76412 59890 76468 59892
rect 76412 59838 76414 59890
rect 76414 59838 76466 59890
rect 76466 59838 76468 59890
rect 76412 59836 76468 59838
rect 78092 59948 78148 60004
rect 77308 59778 77364 59780
rect 77308 59726 77310 59778
rect 77310 59726 77362 59778
rect 77362 59726 77364 59778
rect 77308 59724 77364 59726
rect 77532 59612 77588 59668
rect 76972 58940 77028 58996
rect 77084 58268 77140 58324
rect 76524 58210 76580 58212
rect 76524 58158 76526 58210
rect 76526 58158 76578 58210
rect 76578 58158 76580 58210
rect 76524 58156 76580 58158
rect 76972 57820 77028 57876
rect 76860 57762 76916 57764
rect 76860 57710 76862 57762
rect 76862 57710 76914 57762
rect 76914 57710 76916 57762
rect 76860 57708 76916 57710
rect 77084 57708 77140 57764
rect 77196 58156 77252 58212
rect 76524 57596 76580 57652
rect 75404 56588 75460 56644
rect 75852 56140 75908 56196
rect 75740 56082 75796 56084
rect 75740 56030 75742 56082
rect 75742 56030 75794 56082
rect 75794 56030 75796 56082
rect 75740 56028 75796 56030
rect 75852 55468 75908 55524
rect 75740 55356 75796 55412
rect 75404 53900 75460 53956
rect 75292 53170 75348 53172
rect 75292 53118 75294 53170
rect 75294 53118 75346 53170
rect 75346 53118 75348 53170
rect 75292 53116 75348 53118
rect 75852 54572 75908 54628
rect 75740 52892 75796 52948
rect 74620 50540 74676 50596
rect 74956 51996 75012 52052
rect 75068 51548 75124 51604
rect 75068 51100 75124 51156
rect 74956 50428 75012 50484
rect 74284 48412 74340 48468
rect 75180 50370 75236 50372
rect 75180 50318 75182 50370
rect 75182 50318 75234 50370
rect 75234 50318 75236 50370
rect 75180 50316 75236 50318
rect 74396 44434 74452 44436
rect 74396 44382 74398 44434
rect 74398 44382 74450 44434
rect 74450 44382 74452 44434
rect 74396 44380 74452 44382
rect 72716 41132 72772 41188
rect 71596 36370 71652 36372
rect 71596 36318 71598 36370
rect 71598 36318 71650 36370
rect 71650 36318 71652 36370
rect 71596 36316 71652 36318
rect 73388 36876 73444 36932
rect 74060 41356 74116 41412
rect 73948 40460 74004 40516
rect 73836 39676 73892 39732
rect 75068 49532 75124 49588
rect 75180 50092 75236 50148
rect 75180 49084 75236 49140
rect 74732 47292 74788 47348
rect 75068 46786 75124 46788
rect 75068 46734 75070 46786
rect 75070 46734 75122 46786
rect 75122 46734 75124 46786
rect 75068 46732 75124 46734
rect 75516 51884 75572 51940
rect 75852 50594 75908 50596
rect 75852 50542 75854 50594
rect 75854 50542 75906 50594
rect 75906 50542 75908 50594
rect 75852 50540 75908 50542
rect 75964 50092 76020 50148
rect 75628 49980 75684 50036
rect 75516 49922 75572 49924
rect 75516 49870 75518 49922
rect 75518 49870 75570 49922
rect 75570 49870 75572 49922
rect 75516 49868 75572 49870
rect 75404 48802 75460 48804
rect 75404 48750 75406 48802
rect 75406 48750 75458 48802
rect 75458 48750 75460 48802
rect 75404 48748 75460 48750
rect 75404 48524 75460 48580
rect 75068 44604 75124 44660
rect 75180 42530 75236 42532
rect 75180 42478 75182 42530
rect 75182 42478 75234 42530
rect 75234 42478 75236 42530
rect 75180 42476 75236 42478
rect 74620 41132 74676 41188
rect 75292 41692 75348 41748
rect 75292 41132 75348 41188
rect 74732 41020 74788 41076
rect 75292 40962 75348 40964
rect 75292 40910 75294 40962
rect 75294 40910 75346 40962
rect 75346 40910 75348 40962
rect 75292 40908 75348 40910
rect 74844 39730 74900 39732
rect 74844 39678 74846 39730
rect 74846 39678 74898 39730
rect 74898 39678 74900 39730
rect 74844 39676 74900 39678
rect 75180 39676 75236 39732
rect 74844 38946 74900 38948
rect 74844 38894 74846 38946
rect 74846 38894 74898 38946
rect 74898 38894 74900 38946
rect 74844 38892 74900 38894
rect 74956 38780 75012 38836
rect 76300 56476 76356 56532
rect 76188 56028 76244 56084
rect 76412 56028 76468 56084
rect 78204 59724 78260 59780
rect 78876 61964 78932 62020
rect 79324 64146 79380 64148
rect 79324 64094 79326 64146
rect 79326 64094 79378 64146
rect 79378 64094 79380 64146
rect 79324 64092 79380 64094
rect 79212 63196 79268 63252
rect 79324 63308 79380 63364
rect 79100 62412 79156 62468
rect 78988 61404 79044 61460
rect 78876 60956 78932 61012
rect 78764 60786 78820 60788
rect 78764 60734 78766 60786
rect 78766 60734 78818 60786
rect 78818 60734 78820 60786
rect 78764 60732 78820 60734
rect 78428 59836 78484 59892
rect 78204 58492 78260 58548
rect 78316 58716 78372 58772
rect 77644 58322 77700 58324
rect 77644 58270 77646 58322
rect 77646 58270 77698 58322
rect 77698 58270 77700 58322
rect 77644 58268 77700 58270
rect 78204 58322 78260 58324
rect 78204 58270 78206 58322
rect 78206 58270 78258 58322
rect 78258 58270 78260 58322
rect 78204 58268 78260 58270
rect 77420 58044 77476 58100
rect 77308 57036 77364 57092
rect 77420 57148 77476 57204
rect 77196 56364 77252 56420
rect 76524 55356 76580 55412
rect 76524 55186 76580 55188
rect 76524 55134 76526 55186
rect 76526 55134 76578 55186
rect 76578 55134 76580 55186
rect 76524 55132 76580 55134
rect 76188 54572 76244 54628
rect 76412 54626 76468 54628
rect 76412 54574 76414 54626
rect 76414 54574 76466 54626
rect 76466 54574 76468 54626
rect 76412 54572 76468 54574
rect 77084 56082 77140 56084
rect 77084 56030 77086 56082
rect 77086 56030 77138 56082
rect 77138 56030 77140 56082
rect 77084 56028 77140 56030
rect 76748 54626 76804 54628
rect 76748 54574 76750 54626
rect 76750 54574 76802 54626
rect 76802 54574 76804 54626
rect 76748 54572 76804 54574
rect 76412 53676 76468 53732
rect 76636 53618 76692 53620
rect 76636 53566 76638 53618
rect 76638 53566 76690 53618
rect 76690 53566 76692 53618
rect 76636 53564 76692 53566
rect 76748 52892 76804 52948
rect 76860 52220 76916 52276
rect 76188 50204 76244 50260
rect 76412 50034 76468 50036
rect 76412 49982 76414 50034
rect 76414 49982 76466 50034
rect 76466 49982 76468 50034
rect 76412 49980 76468 49982
rect 76188 49138 76244 49140
rect 76188 49086 76190 49138
rect 76190 49086 76242 49138
rect 76242 49086 76244 49138
rect 76188 49084 76244 49086
rect 75852 46898 75908 46900
rect 75852 46846 75854 46898
rect 75854 46846 75906 46898
rect 75906 46846 75908 46898
rect 75852 46844 75908 46846
rect 75516 46786 75572 46788
rect 75516 46734 75518 46786
rect 75518 46734 75570 46786
rect 75570 46734 75572 46786
rect 75516 46732 75572 46734
rect 76748 50316 76804 50372
rect 76860 50428 76916 50484
rect 77196 55186 77252 55188
rect 77196 55134 77198 55186
rect 77198 55134 77250 55186
rect 77250 55134 77252 55186
rect 77196 55132 77252 55134
rect 77420 56588 77476 56644
rect 78428 58492 78484 58548
rect 78988 59330 79044 59332
rect 78988 59278 78990 59330
rect 78990 59278 79042 59330
rect 79042 59278 79044 59330
rect 78988 59276 79044 59278
rect 78540 58210 78596 58212
rect 78540 58158 78542 58210
rect 78542 58158 78594 58210
rect 78594 58158 78596 58210
rect 78540 58156 78596 58158
rect 79660 64092 79716 64148
rect 79660 63644 79716 63700
rect 80108 65324 80164 65380
rect 79996 64706 80052 64708
rect 79996 64654 79998 64706
rect 79998 64654 80050 64706
rect 80050 64654 80052 64706
rect 79996 64652 80052 64654
rect 79884 64204 79940 64260
rect 79996 63980 80052 64036
rect 79548 62860 79604 62916
rect 79884 63756 79940 63812
rect 79436 62466 79492 62468
rect 79436 62414 79438 62466
rect 79438 62414 79490 62466
rect 79490 62414 79492 62466
rect 79436 62412 79492 62414
rect 79772 62188 79828 62244
rect 79660 61964 79716 62020
rect 79436 61292 79492 61348
rect 79324 60898 79380 60900
rect 79324 60846 79326 60898
rect 79326 60846 79378 60898
rect 79378 60846 79380 60898
rect 79324 60844 79380 60846
rect 79660 61346 79716 61348
rect 79660 61294 79662 61346
rect 79662 61294 79714 61346
rect 79714 61294 79716 61346
rect 79660 61292 79716 61294
rect 79660 60956 79716 61012
rect 79100 58380 79156 58436
rect 78876 58044 78932 58100
rect 78428 57820 78484 57876
rect 78540 57932 78596 57988
rect 78876 57874 78932 57876
rect 78876 57822 78878 57874
rect 78878 57822 78930 57874
rect 78930 57822 78932 57874
rect 78876 57820 78932 57822
rect 78316 57148 78372 57204
rect 78988 56978 79044 56980
rect 78988 56926 78990 56978
rect 78990 56926 79042 56978
rect 79042 56926 79044 56978
rect 78988 56924 79044 56926
rect 77756 56252 77812 56308
rect 77868 56476 77924 56532
rect 78428 55804 78484 55860
rect 78204 55244 78260 55300
rect 77644 54684 77700 54740
rect 77756 54514 77812 54516
rect 77756 54462 77758 54514
rect 77758 54462 77810 54514
rect 77810 54462 77812 54514
rect 77756 54460 77812 54462
rect 77308 53116 77364 53172
rect 77084 51378 77140 51380
rect 77084 51326 77086 51378
rect 77086 51326 77138 51378
rect 77138 51326 77140 51378
rect 77084 51324 77140 51326
rect 77420 51884 77476 51940
rect 77084 50316 77140 50372
rect 77196 50482 77252 50484
rect 77196 50430 77198 50482
rect 77198 50430 77250 50482
rect 77250 50430 77252 50482
rect 77196 50428 77252 50430
rect 76524 48636 76580 48692
rect 76524 48412 76580 48468
rect 76412 47404 76468 47460
rect 76300 46844 76356 46900
rect 76748 48242 76804 48244
rect 76748 48190 76750 48242
rect 76750 48190 76802 48242
rect 76802 48190 76804 48242
rect 76748 48188 76804 48190
rect 76076 46002 76132 46004
rect 76076 45950 76078 46002
rect 76078 45950 76130 46002
rect 76130 45950 76132 46002
rect 76076 45948 76132 45950
rect 76076 44604 76132 44660
rect 75628 44380 75684 44436
rect 75964 44380 76020 44436
rect 75740 42754 75796 42756
rect 75740 42702 75742 42754
rect 75742 42702 75794 42754
rect 75794 42702 75796 42754
rect 75740 42700 75796 42702
rect 75852 41298 75908 41300
rect 75852 41246 75854 41298
rect 75854 41246 75906 41298
rect 75906 41246 75908 41298
rect 75852 41244 75908 41246
rect 75404 39618 75460 39620
rect 75404 39566 75406 39618
rect 75406 39566 75458 39618
rect 75458 39566 75460 39618
rect 75404 39564 75460 39566
rect 74060 36876 74116 36932
rect 71148 34300 71204 34356
rect 70812 33292 70868 33348
rect 70252 33068 70308 33124
rect 69580 32450 69636 32452
rect 69580 32398 69582 32450
rect 69582 32398 69634 32450
rect 69634 32398 69636 32450
rect 69580 32396 69636 32398
rect 69244 32338 69300 32340
rect 69244 32286 69246 32338
rect 69246 32286 69298 32338
rect 69298 32286 69300 32338
rect 69244 32284 69300 32286
rect 70364 33180 70420 33236
rect 71372 33180 71428 33236
rect 70924 32562 70980 32564
rect 70924 32510 70926 32562
rect 70926 32510 70978 32562
rect 70978 32510 70980 32562
rect 70924 32508 70980 32510
rect 69356 31724 69412 31780
rect 67676 31666 67732 31668
rect 67676 31614 67678 31666
rect 67678 31614 67730 31666
rect 67730 31614 67732 31666
rect 67676 31612 67732 31614
rect 56140 3388 56196 3444
rect 54348 3276 54404 3332
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 45276 2716 45332 2772
rect 56700 3442 56756 3444
rect 56700 3390 56702 3442
rect 56702 3390 56754 3442
rect 56754 3390 56756 3442
rect 56700 3388 56756 3390
rect 57036 2940 57092 2996
rect 72380 34972 72436 35028
rect 72156 34914 72212 34916
rect 72156 34862 72158 34914
rect 72158 34862 72210 34914
rect 72210 34862 72212 34914
rect 72156 34860 72212 34862
rect 72604 34860 72660 34916
rect 72044 34636 72100 34692
rect 72604 34076 72660 34132
rect 73052 33122 73108 33124
rect 73052 33070 73054 33122
rect 73054 33070 73106 33122
rect 73106 33070 73108 33122
rect 73052 33068 73108 33070
rect 72604 32786 72660 32788
rect 72604 32734 72606 32786
rect 72606 32734 72658 32786
rect 72658 32734 72660 32786
rect 72604 32732 72660 32734
rect 73276 32562 73332 32564
rect 73276 32510 73278 32562
rect 73278 32510 73330 32562
rect 73330 32510 73332 32562
rect 73276 32508 73332 32510
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 67788 3442 67844 3444
rect 67788 3390 67790 3442
rect 67790 3390 67842 3442
rect 67842 3390 67844 3442
rect 67788 3388 67844 3390
rect 68796 3442 68852 3444
rect 68796 3390 68798 3442
rect 68798 3390 68850 3442
rect 68850 3390 68852 3442
rect 68796 3388 68852 3390
rect 57372 2828 57428 2884
rect 73500 34972 73556 35028
rect 73724 34914 73780 34916
rect 73724 34862 73726 34914
rect 73726 34862 73778 34914
rect 73778 34862 73780 34914
rect 73724 34860 73780 34862
rect 74620 36876 74676 36932
rect 75516 40460 75572 40516
rect 75628 38668 75684 38724
rect 75852 38050 75908 38052
rect 75852 37998 75854 38050
rect 75854 37998 75906 38050
rect 75906 37998 75908 38050
rect 75852 37996 75908 37998
rect 75964 37938 76020 37940
rect 75964 37886 75966 37938
rect 75966 37886 76018 37938
rect 76018 37886 76020 37938
rect 75964 37884 76020 37886
rect 75852 37378 75908 37380
rect 75852 37326 75854 37378
rect 75854 37326 75906 37378
rect 75906 37326 75908 37378
rect 75852 37324 75908 37326
rect 75404 36876 75460 36932
rect 74284 35868 74340 35924
rect 74620 36428 74676 36484
rect 74396 35756 74452 35812
rect 73500 34354 73556 34356
rect 73500 34302 73502 34354
rect 73502 34302 73554 34354
rect 73554 34302 73556 34354
rect 73500 34300 73556 34302
rect 73836 34130 73892 34132
rect 73836 34078 73838 34130
rect 73838 34078 73890 34130
rect 73890 34078 73892 34130
rect 73836 34076 73892 34078
rect 74956 36482 75012 36484
rect 74956 36430 74958 36482
rect 74958 36430 75010 36482
rect 75010 36430 75012 36482
rect 74956 36428 75012 36430
rect 76524 44434 76580 44436
rect 76524 44382 76526 44434
rect 76526 44382 76578 44434
rect 76578 44382 76580 44434
rect 76524 44380 76580 44382
rect 76748 42924 76804 42980
rect 76188 42530 76244 42532
rect 76188 42478 76190 42530
rect 76190 42478 76242 42530
rect 76242 42478 76244 42530
rect 76188 42476 76244 42478
rect 78092 53618 78148 53620
rect 78092 53566 78094 53618
rect 78094 53566 78146 53618
rect 78146 53566 78148 53618
rect 78092 53564 78148 53566
rect 78876 55858 78932 55860
rect 78876 55806 78878 55858
rect 78878 55806 78930 55858
rect 78930 55806 78932 55858
rect 78876 55804 78932 55806
rect 79324 59218 79380 59220
rect 79324 59166 79326 59218
rect 79326 59166 79378 59218
rect 79378 59166 79380 59218
rect 79324 59164 79380 59166
rect 79324 58044 79380 58100
rect 79324 57708 79380 57764
rect 79436 58156 79492 58212
rect 80332 64988 80388 65044
rect 80220 64092 80276 64148
rect 80444 63868 80500 63924
rect 80332 62412 80388 62468
rect 80108 61964 80164 62020
rect 79772 60060 79828 60116
rect 79996 60396 80052 60452
rect 80220 61852 80276 61908
rect 80780 66332 80836 66388
rect 81564 67058 81620 67060
rect 81564 67006 81566 67058
rect 81566 67006 81618 67058
rect 81618 67006 81620 67058
rect 81564 67004 81620 67006
rect 81004 65772 81060 65828
rect 80892 65660 80948 65716
rect 81004 65548 81060 65604
rect 81276 65882 81332 65884
rect 81276 65830 81278 65882
rect 81278 65830 81330 65882
rect 81330 65830 81332 65882
rect 81276 65828 81332 65830
rect 81380 65882 81436 65884
rect 81380 65830 81382 65882
rect 81382 65830 81434 65882
rect 81434 65830 81436 65882
rect 81380 65828 81436 65830
rect 81484 65882 81540 65884
rect 81484 65830 81486 65882
rect 81486 65830 81538 65882
rect 81538 65830 81540 65882
rect 81484 65828 81540 65830
rect 81116 65324 81172 65380
rect 81228 64988 81284 65044
rect 81004 64540 81060 64596
rect 80556 62524 80612 62580
rect 80668 63196 80724 63252
rect 80668 62860 80724 62916
rect 80780 62188 80836 62244
rect 81276 64314 81332 64316
rect 81276 64262 81278 64314
rect 81278 64262 81330 64314
rect 81330 64262 81332 64314
rect 81276 64260 81332 64262
rect 81380 64314 81436 64316
rect 81380 64262 81382 64314
rect 81382 64262 81434 64314
rect 81434 64262 81436 64314
rect 81380 64260 81436 64262
rect 81484 64314 81540 64316
rect 81484 64262 81486 64314
rect 81486 64262 81538 64314
rect 81538 64262 81540 64314
rect 81484 64260 81540 64262
rect 81116 64092 81172 64148
rect 81564 63922 81620 63924
rect 81564 63870 81566 63922
rect 81566 63870 81618 63922
rect 81618 63870 81620 63922
rect 81564 63868 81620 63870
rect 81900 70140 81956 70196
rect 81900 69468 81956 69524
rect 82124 69298 82180 69300
rect 82124 69246 82126 69298
rect 82126 69246 82178 69298
rect 82178 69246 82180 69298
rect 82124 69244 82180 69246
rect 82908 70476 82964 70532
rect 83020 70700 83076 70756
rect 82684 69244 82740 69300
rect 83356 70476 83412 70532
rect 82572 68908 82628 68964
rect 82572 67842 82628 67844
rect 82572 67790 82574 67842
rect 82574 67790 82626 67842
rect 82626 67790 82628 67842
rect 82572 67788 82628 67790
rect 82572 67116 82628 67172
rect 82012 66780 82068 66836
rect 81900 66444 81956 66500
rect 82124 66444 82180 66500
rect 81900 65548 81956 65604
rect 81788 64540 81844 64596
rect 82348 66386 82404 66388
rect 82348 66334 82350 66386
rect 82350 66334 82402 66386
rect 82402 66334 82404 66386
rect 82348 66332 82404 66334
rect 82236 65100 82292 65156
rect 82012 64146 82068 64148
rect 82012 64094 82014 64146
rect 82014 64094 82066 64146
rect 82066 64094 82068 64146
rect 82012 64092 82068 64094
rect 81788 63922 81844 63924
rect 81788 63870 81790 63922
rect 81790 63870 81842 63922
rect 81842 63870 81844 63922
rect 81788 63868 81844 63870
rect 81564 63196 81620 63252
rect 81004 62972 81060 63028
rect 82348 63308 82404 63364
rect 82460 64204 82516 64260
rect 81276 62746 81332 62748
rect 81276 62694 81278 62746
rect 81278 62694 81330 62746
rect 81330 62694 81332 62746
rect 81276 62692 81332 62694
rect 81380 62746 81436 62748
rect 81380 62694 81382 62746
rect 81382 62694 81434 62746
rect 81434 62694 81436 62746
rect 81380 62692 81436 62694
rect 81484 62746 81540 62748
rect 81484 62694 81486 62746
rect 81486 62694 81538 62746
rect 81538 62694 81540 62746
rect 81484 62692 81540 62694
rect 81900 62524 81956 62580
rect 81340 62466 81396 62468
rect 81340 62414 81342 62466
rect 81342 62414 81394 62466
rect 81394 62414 81396 62466
rect 81340 62412 81396 62414
rect 81676 62354 81732 62356
rect 81676 62302 81678 62354
rect 81678 62302 81730 62354
rect 81730 62302 81732 62354
rect 81676 62300 81732 62302
rect 82124 62300 82180 62356
rect 80220 60508 80276 60564
rect 80220 59836 80276 59892
rect 80892 59388 80948 59444
rect 79996 59164 80052 59220
rect 79772 59106 79828 59108
rect 79772 59054 79774 59106
rect 79774 59054 79826 59106
rect 79826 59054 79828 59106
rect 79772 59052 79828 59054
rect 79772 58434 79828 58436
rect 79772 58382 79774 58434
rect 79774 58382 79826 58434
rect 79826 58382 79828 58434
rect 79772 58380 79828 58382
rect 79548 57762 79604 57764
rect 79548 57710 79550 57762
rect 79550 57710 79602 57762
rect 79602 57710 79604 57762
rect 79548 57708 79604 57710
rect 79548 56924 79604 56980
rect 79436 56588 79492 56644
rect 79100 54572 79156 54628
rect 79212 54348 79268 54404
rect 79548 54572 79604 54628
rect 78764 53676 78820 53732
rect 77644 53170 77700 53172
rect 77644 53118 77646 53170
rect 77646 53118 77698 53170
rect 77698 53118 77700 53170
rect 77644 53116 77700 53118
rect 77644 52274 77700 52276
rect 77644 52222 77646 52274
rect 77646 52222 77698 52274
rect 77698 52222 77700 52274
rect 77644 52220 77700 52222
rect 78428 53170 78484 53172
rect 78428 53118 78430 53170
rect 78430 53118 78482 53170
rect 78482 53118 78484 53170
rect 78428 53116 78484 53118
rect 77308 49026 77364 49028
rect 77308 48974 77310 49026
rect 77310 48974 77362 49026
rect 77362 48974 77364 49026
rect 77308 48972 77364 48974
rect 77644 50316 77700 50372
rect 77756 48972 77812 49028
rect 77532 48188 77588 48244
rect 77644 48636 77700 48692
rect 77644 47516 77700 47572
rect 77196 47458 77252 47460
rect 77196 47406 77198 47458
rect 77198 47406 77250 47458
rect 77250 47406 77252 47458
rect 77196 47404 77252 47406
rect 77420 45724 77476 45780
rect 77084 43596 77140 43652
rect 77196 45052 77252 45108
rect 78316 52946 78372 52948
rect 78316 52894 78318 52946
rect 78318 52894 78370 52946
rect 78370 52894 78372 52946
rect 78316 52892 78372 52894
rect 79100 52946 79156 52948
rect 79100 52894 79102 52946
rect 79102 52894 79154 52946
rect 79154 52894 79156 52946
rect 79100 52892 79156 52894
rect 78764 52556 78820 52612
rect 79100 52556 79156 52612
rect 78316 51490 78372 51492
rect 78316 51438 78318 51490
rect 78318 51438 78370 51490
rect 78370 51438 78372 51490
rect 78316 51436 78372 51438
rect 78204 51378 78260 51380
rect 78204 51326 78206 51378
rect 78206 51326 78258 51378
rect 78258 51326 78260 51378
rect 78204 51324 78260 51326
rect 79436 51490 79492 51492
rect 79436 51438 79438 51490
rect 79438 51438 79490 51490
rect 79490 51438 79492 51490
rect 79436 51436 79492 51438
rect 79100 50204 79156 50260
rect 78764 50092 78820 50148
rect 78428 49868 78484 49924
rect 77980 49084 78036 49140
rect 78428 49084 78484 49140
rect 78652 48972 78708 49028
rect 78092 48412 78148 48468
rect 78316 48466 78372 48468
rect 78316 48414 78318 48466
rect 78318 48414 78370 48466
rect 78370 48414 78372 48466
rect 78316 48412 78372 48414
rect 78652 48188 78708 48244
rect 78092 48076 78148 48132
rect 79548 50594 79604 50596
rect 79548 50542 79550 50594
rect 79550 50542 79602 50594
rect 79602 50542 79604 50594
rect 79548 50540 79604 50542
rect 81676 62076 81732 62132
rect 81452 61740 81508 61796
rect 81276 61178 81332 61180
rect 81276 61126 81278 61178
rect 81278 61126 81330 61178
rect 81330 61126 81332 61178
rect 81276 61124 81332 61126
rect 81380 61178 81436 61180
rect 81380 61126 81382 61178
rect 81382 61126 81434 61178
rect 81434 61126 81436 61178
rect 81380 61124 81436 61126
rect 81484 61178 81540 61180
rect 81484 61126 81486 61178
rect 81486 61126 81538 61178
rect 81538 61126 81540 61178
rect 81484 61124 81540 61126
rect 81676 60844 81732 60900
rect 82236 62636 82292 62692
rect 82460 62412 82516 62468
rect 82236 61682 82292 61684
rect 82236 61630 82238 61682
rect 82238 61630 82290 61682
rect 82290 61630 82292 61682
rect 82236 61628 82292 61630
rect 82348 60898 82404 60900
rect 82348 60846 82350 60898
rect 82350 60846 82402 60898
rect 82402 60846 82404 60898
rect 82348 60844 82404 60846
rect 81452 60396 81508 60452
rect 81340 60172 81396 60228
rect 81676 60002 81732 60004
rect 81676 59950 81678 60002
rect 81678 59950 81730 60002
rect 81730 59950 81732 60002
rect 81676 59948 81732 59950
rect 81116 59724 81172 59780
rect 82236 60508 82292 60564
rect 81900 59724 81956 59780
rect 82012 59948 82068 60004
rect 81276 59610 81332 59612
rect 81276 59558 81278 59610
rect 81278 59558 81330 59610
rect 81330 59558 81332 59610
rect 81276 59556 81332 59558
rect 81380 59610 81436 59612
rect 81380 59558 81382 59610
rect 81382 59558 81434 59610
rect 81434 59558 81436 59610
rect 81380 59556 81436 59558
rect 81484 59610 81540 59612
rect 81484 59558 81486 59610
rect 81486 59558 81538 59610
rect 81538 59558 81540 59610
rect 81484 59556 81540 59558
rect 81004 58716 81060 58772
rect 80220 58546 80276 58548
rect 80220 58494 80222 58546
rect 80222 58494 80274 58546
rect 80274 58494 80276 58546
rect 80220 58492 80276 58494
rect 81564 58322 81620 58324
rect 81564 58270 81566 58322
rect 81566 58270 81618 58322
rect 81618 58270 81620 58322
rect 81564 58268 81620 58270
rect 82124 59500 82180 59556
rect 82236 59052 82292 59108
rect 82124 58940 82180 58996
rect 81676 58156 81732 58212
rect 80668 57932 80724 57988
rect 81276 58042 81332 58044
rect 81276 57990 81278 58042
rect 81278 57990 81330 58042
rect 81330 57990 81332 58042
rect 81276 57988 81332 57990
rect 81380 58042 81436 58044
rect 81380 57990 81382 58042
rect 81382 57990 81434 58042
rect 81434 57990 81436 58042
rect 81380 57988 81436 57990
rect 81484 58042 81540 58044
rect 81484 57990 81486 58042
rect 81486 57990 81538 58042
rect 81538 57990 81540 58042
rect 81484 57988 81540 57990
rect 80332 57820 80388 57876
rect 82012 57874 82068 57876
rect 82012 57822 82014 57874
rect 82014 57822 82066 57874
rect 82066 57822 82068 57874
rect 82012 57820 82068 57822
rect 79996 57036 80052 57092
rect 80668 57762 80724 57764
rect 80668 57710 80670 57762
rect 80670 57710 80722 57762
rect 80722 57710 80724 57762
rect 80668 57708 80724 57710
rect 81340 57762 81396 57764
rect 81340 57710 81342 57762
rect 81342 57710 81394 57762
rect 81394 57710 81396 57762
rect 81340 57708 81396 57710
rect 80556 56924 80612 56980
rect 81116 56978 81172 56980
rect 81116 56926 81118 56978
rect 81118 56926 81170 56978
rect 81170 56926 81172 56978
rect 81116 56924 81172 56926
rect 80556 56588 80612 56644
rect 80332 56306 80388 56308
rect 80332 56254 80334 56306
rect 80334 56254 80386 56306
rect 80386 56254 80388 56306
rect 80332 56252 80388 56254
rect 79772 55298 79828 55300
rect 79772 55246 79774 55298
rect 79774 55246 79826 55298
rect 79826 55246 79828 55298
rect 79772 55244 79828 55246
rect 79996 51490 80052 51492
rect 79996 51438 79998 51490
rect 79998 51438 80050 51490
rect 80050 51438 80052 51490
rect 79996 51436 80052 51438
rect 79884 51378 79940 51380
rect 79884 51326 79886 51378
rect 79886 51326 79938 51378
rect 79938 51326 79940 51378
rect 79884 51324 79940 51326
rect 79212 49644 79268 49700
rect 79100 49026 79156 49028
rect 79100 48974 79102 49026
rect 79102 48974 79154 49026
rect 79154 48974 79156 49026
rect 79100 48972 79156 48974
rect 79100 45778 79156 45780
rect 79100 45726 79102 45778
rect 79102 45726 79154 45778
rect 79154 45726 79156 45778
rect 79100 45724 79156 45726
rect 77868 45612 77924 45668
rect 77756 45106 77812 45108
rect 77756 45054 77758 45106
rect 77758 45054 77810 45106
rect 77810 45054 77812 45106
rect 77756 45052 77812 45054
rect 77756 44434 77812 44436
rect 77756 44382 77758 44434
rect 77758 44382 77810 44434
rect 77810 44382 77812 44434
rect 77756 44380 77812 44382
rect 79212 45612 79268 45668
rect 78540 44210 78596 44212
rect 78540 44158 78542 44210
rect 78542 44158 78594 44210
rect 78594 44158 78596 44210
rect 78540 44156 78596 44158
rect 77756 43708 77812 43764
rect 77420 42978 77476 42980
rect 77420 42926 77422 42978
rect 77422 42926 77474 42978
rect 77474 42926 77476 42978
rect 77420 42924 77476 42926
rect 77868 43650 77924 43652
rect 77868 43598 77870 43650
rect 77870 43598 77922 43650
rect 77922 43598 77924 43650
rect 77868 43596 77924 43598
rect 81788 56754 81844 56756
rect 81788 56702 81790 56754
rect 81790 56702 81842 56754
rect 81842 56702 81844 56754
rect 81788 56700 81844 56702
rect 81452 56588 81508 56644
rect 81900 56588 81956 56644
rect 81276 56474 81332 56476
rect 81276 56422 81278 56474
rect 81278 56422 81330 56474
rect 81330 56422 81332 56474
rect 81276 56420 81332 56422
rect 81380 56474 81436 56476
rect 81380 56422 81382 56474
rect 81382 56422 81434 56474
rect 81434 56422 81436 56474
rect 81380 56420 81436 56422
rect 81484 56474 81540 56476
rect 81484 56422 81486 56474
rect 81486 56422 81538 56474
rect 81538 56422 81540 56474
rect 81484 56420 81540 56422
rect 81900 56252 81956 56308
rect 81788 55244 81844 55300
rect 81276 54906 81332 54908
rect 81276 54854 81278 54906
rect 81278 54854 81330 54906
rect 81330 54854 81332 54906
rect 81276 54852 81332 54854
rect 81380 54906 81436 54908
rect 81380 54854 81382 54906
rect 81382 54854 81434 54906
rect 81434 54854 81436 54906
rect 81380 54852 81436 54854
rect 81484 54906 81540 54908
rect 81484 54854 81486 54906
rect 81486 54854 81538 54906
rect 81538 54854 81540 54906
rect 81484 54852 81540 54854
rect 80668 54460 80724 54516
rect 80556 54402 80612 54404
rect 80556 54350 80558 54402
rect 80558 54350 80610 54402
rect 80610 54350 80612 54402
rect 80556 54348 80612 54350
rect 80220 53116 80276 53172
rect 82124 55244 82180 55300
rect 81276 53338 81332 53340
rect 81276 53286 81278 53338
rect 81278 53286 81330 53338
rect 81330 53286 81332 53338
rect 81276 53284 81332 53286
rect 81380 53338 81436 53340
rect 81380 53286 81382 53338
rect 81382 53286 81434 53338
rect 81434 53286 81436 53338
rect 81380 53284 81436 53286
rect 81484 53338 81540 53340
rect 81484 53286 81486 53338
rect 81486 53286 81538 53338
rect 81538 53286 81540 53338
rect 81484 53284 81540 53286
rect 81276 51770 81332 51772
rect 81276 51718 81278 51770
rect 81278 51718 81330 51770
rect 81330 51718 81332 51770
rect 81276 51716 81332 51718
rect 81380 51770 81436 51772
rect 81380 51718 81382 51770
rect 81382 51718 81434 51770
rect 81434 51718 81436 51770
rect 81380 51716 81436 51718
rect 81484 51770 81540 51772
rect 81484 51718 81486 51770
rect 81486 51718 81538 51770
rect 81538 51718 81540 51770
rect 81484 51716 81540 51718
rect 82796 65660 82852 65716
rect 82684 65100 82740 65156
rect 83020 68572 83076 68628
rect 83020 67842 83076 67844
rect 83020 67790 83022 67842
rect 83022 67790 83074 67842
rect 83074 67790 83076 67842
rect 83020 67788 83076 67790
rect 83692 70476 83748 70532
rect 83580 69186 83636 69188
rect 83580 69134 83582 69186
rect 83582 69134 83634 69186
rect 83634 69134 83636 69186
rect 83580 69132 83636 69134
rect 83468 68908 83524 68964
rect 83244 67170 83300 67172
rect 83244 67118 83246 67170
rect 83246 67118 83298 67170
rect 83298 67118 83300 67170
rect 83244 67116 83300 67118
rect 83132 67058 83188 67060
rect 83132 67006 83134 67058
rect 83134 67006 83186 67058
rect 83186 67006 83188 67058
rect 83132 67004 83188 67006
rect 83244 66108 83300 66164
rect 83692 67788 83748 67844
rect 83580 67004 83636 67060
rect 83580 66050 83636 66052
rect 83580 65998 83582 66050
rect 83582 65998 83634 66050
rect 83634 65998 83636 66050
rect 83580 65996 83636 65998
rect 82908 64988 82964 65044
rect 83020 65212 83076 65268
rect 82684 64652 82740 64708
rect 82796 64316 82852 64372
rect 82908 64146 82964 64148
rect 82908 64094 82910 64146
rect 82910 64094 82962 64146
rect 82962 64094 82964 64146
rect 82908 64092 82964 64094
rect 83580 64876 83636 64932
rect 83132 64764 83188 64820
rect 83244 64706 83300 64708
rect 83244 64654 83246 64706
rect 83246 64654 83298 64706
rect 83298 64654 83300 64706
rect 83244 64652 83300 64654
rect 82796 63868 82852 63924
rect 82908 63756 82964 63812
rect 82684 62636 82740 62692
rect 82796 63644 82852 63700
rect 82796 62076 82852 62132
rect 82796 60898 82852 60900
rect 82796 60846 82798 60898
rect 82798 60846 82850 60898
rect 82850 60846 82852 60898
rect 82796 60844 82852 60846
rect 82572 59106 82628 59108
rect 82572 59054 82574 59106
rect 82574 59054 82626 59106
rect 82626 59054 82628 59106
rect 82572 59052 82628 59054
rect 82348 56700 82404 56756
rect 82348 52444 82404 52500
rect 83132 63644 83188 63700
rect 83020 63138 83076 63140
rect 83020 63086 83022 63138
rect 83022 63086 83074 63138
rect 83074 63086 83076 63138
rect 83020 63084 83076 63086
rect 83020 62860 83076 62916
rect 83244 62524 83300 62580
rect 83244 62354 83300 62356
rect 83244 62302 83246 62354
rect 83246 62302 83298 62354
rect 83298 62302 83300 62354
rect 83244 62300 83300 62302
rect 83580 63868 83636 63924
rect 84028 74844 84084 74900
rect 83916 72268 83972 72324
rect 83916 68572 83972 68628
rect 83916 67228 83972 67284
rect 83804 67116 83860 67172
rect 84588 75516 84644 75572
rect 85260 75628 85316 75684
rect 86044 80498 86100 80500
rect 86044 80446 86046 80498
rect 86046 80446 86098 80498
rect 86098 80446 86100 80498
rect 86044 80444 86100 80446
rect 86268 79714 86324 79716
rect 86268 79662 86270 79714
rect 86270 79662 86322 79714
rect 86322 79662 86324 79714
rect 86268 79660 86324 79662
rect 86044 79602 86100 79604
rect 86044 79550 86046 79602
rect 86046 79550 86098 79602
rect 86098 79550 86100 79602
rect 86044 79548 86100 79550
rect 85932 78764 85988 78820
rect 86156 77196 86212 77252
rect 85708 76636 85764 76692
rect 86044 76860 86100 76916
rect 86044 75740 86100 75796
rect 84476 72322 84532 72324
rect 84476 72270 84478 72322
rect 84478 72270 84530 72322
rect 84530 72270 84532 72322
rect 84476 72268 84532 72270
rect 85372 71820 85428 71876
rect 84252 71148 84308 71204
rect 85708 71202 85764 71204
rect 85708 71150 85710 71202
rect 85710 71150 85762 71202
rect 85762 71150 85764 71202
rect 85708 71148 85764 71150
rect 86380 76354 86436 76356
rect 86380 76302 86382 76354
rect 86382 76302 86434 76354
rect 86434 76302 86436 76354
rect 86380 76300 86436 76302
rect 86716 80668 86772 80724
rect 87724 84418 87780 84420
rect 87724 84366 87726 84418
rect 87726 84366 87778 84418
rect 87778 84366 87780 84418
rect 87724 84364 87780 84366
rect 87612 83298 87668 83300
rect 87612 83246 87614 83298
rect 87614 83246 87666 83298
rect 87666 83246 87668 83298
rect 87612 83244 87668 83246
rect 87612 82572 87668 82628
rect 86828 80444 86884 80500
rect 86828 79772 86884 79828
rect 87388 79660 87444 79716
rect 87724 78876 87780 78932
rect 87500 78818 87556 78820
rect 87500 78766 87502 78818
rect 87502 78766 87554 78818
rect 87554 78766 87556 78818
rect 87500 78764 87556 78766
rect 87612 78034 87668 78036
rect 87612 77982 87614 78034
rect 87614 77982 87666 78034
rect 87666 77982 87668 78034
rect 87612 77980 87668 77982
rect 86716 77084 86772 77140
rect 86716 75794 86772 75796
rect 86716 75742 86718 75794
rect 86718 75742 86770 75794
rect 86770 75742 86772 75794
rect 86716 75740 86772 75742
rect 86380 75682 86436 75684
rect 86380 75630 86382 75682
rect 86382 75630 86434 75682
rect 86434 75630 86436 75682
rect 86380 75628 86436 75630
rect 86604 72492 86660 72548
rect 85932 70866 85988 70868
rect 85932 70814 85934 70866
rect 85934 70814 85986 70866
rect 85986 70814 85988 70866
rect 85932 70812 85988 70814
rect 84588 70754 84644 70756
rect 84588 70702 84590 70754
rect 84590 70702 84642 70754
rect 84642 70702 84644 70754
rect 84588 70700 84644 70702
rect 85372 70082 85428 70084
rect 85372 70030 85374 70082
rect 85374 70030 85426 70082
rect 85426 70030 85428 70082
rect 85372 70028 85428 70030
rect 85596 70028 85652 70084
rect 84364 69468 84420 69524
rect 84476 69410 84532 69412
rect 84476 69358 84478 69410
rect 84478 69358 84530 69410
rect 84530 69358 84532 69410
rect 84476 69356 84532 69358
rect 84364 69186 84420 69188
rect 84364 69134 84366 69186
rect 84366 69134 84418 69186
rect 84418 69134 84420 69186
rect 84364 69132 84420 69134
rect 85260 68908 85316 68964
rect 84252 67842 84308 67844
rect 84252 67790 84254 67842
rect 84254 67790 84306 67842
rect 84306 67790 84308 67842
rect 84252 67788 84308 67790
rect 85148 67676 85204 67732
rect 84252 67340 84308 67396
rect 84700 67340 84756 67396
rect 85260 67564 85316 67620
rect 85372 67282 85428 67284
rect 85372 67230 85374 67282
rect 85374 67230 85426 67282
rect 85426 67230 85428 67282
rect 85372 67228 85428 67230
rect 85484 67170 85540 67172
rect 85484 67118 85486 67170
rect 85486 67118 85538 67170
rect 85538 67118 85540 67170
rect 85484 67116 85540 67118
rect 84028 66332 84084 66388
rect 84252 66162 84308 66164
rect 84252 66110 84254 66162
rect 84254 66110 84306 66162
rect 84306 66110 84308 66162
rect 84252 66108 84308 66110
rect 84140 65996 84196 66052
rect 84364 65660 84420 65716
rect 84140 65548 84196 65604
rect 85372 66220 85428 66276
rect 85372 65772 85428 65828
rect 83916 63922 83972 63924
rect 83916 63870 83918 63922
rect 83918 63870 83970 63922
rect 83970 63870 83972 63922
rect 83916 63868 83972 63870
rect 83804 63026 83860 63028
rect 83804 62974 83806 63026
rect 83806 62974 83858 63026
rect 83858 62974 83860 63026
rect 83804 62972 83860 62974
rect 83916 62914 83972 62916
rect 83916 62862 83918 62914
rect 83918 62862 83970 62914
rect 83970 62862 83972 62914
rect 83916 62860 83972 62862
rect 83580 62412 83636 62468
rect 83692 62354 83748 62356
rect 83692 62302 83694 62354
rect 83694 62302 83746 62354
rect 83746 62302 83748 62354
rect 83692 62300 83748 62302
rect 83468 62188 83524 62244
rect 85484 65996 85540 66052
rect 84812 64034 84868 64036
rect 84812 63982 84814 64034
rect 84814 63982 84866 64034
rect 84866 63982 84868 64034
rect 84812 63980 84868 63982
rect 84924 63868 84980 63924
rect 84364 63196 84420 63252
rect 84028 62412 84084 62468
rect 83916 62300 83972 62356
rect 83468 61570 83524 61572
rect 83468 61518 83470 61570
rect 83470 61518 83522 61570
rect 83522 61518 83524 61570
rect 83468 61516 83524 61518
rect 83244 60786 83300 60788
rect 83244 60734 83246 60786
rect 83246 60734 83298 60786
rect 83298 60734 83300 60786
rect 83244 60732 83300 60734
rect 83692 61628 83748 61684
rect 83580 60284 83636 60340
rect 83132 60114 83188 60116
rect 83132 60062 83134 60114
rect 83134 60062 83186 60114
rect 83186 60062 83188 60114
rect 83132 60060 83188 60062
rect 83468 59442 83524 59444
rect 83468 59390 83470 59442
rect 83470 59390 83522 59442
rect 83522 59390 83524 59442
rect 83468 59388 83524 59390
rect 83132 58604 83188 58660
rect 84476 62972 84532 63028
rect 84364 62578 84420 62580
rect 84364 62526 84366 62578
rect 84366 62526 84418 62578
rect 84418 62526 84420 62578
rect 84364 62524 84420 62526
rect 84364 61346 84420 61348
rect 84364 61294 84366 61346
rect 84366 61294 84418 61346
rect 84418 61294 84420 61346
rect 84364 61292 84420 61294
rect 84252 61068 84308 61124
rect 84140 60898 84196 60900
rect 84140 60846 84142 60898
rect 84142 60846 84194 60898
rect 84194 60846 84196 60898
rect 84140 60844 84196 60846
rect 84252 60786 84308 60788
rect 84252 60734 84254 60786
rect 84254 60734 84306 60786
rect 84306 60734 84308 60786
rect 84252 60732 84308 60734
rect 84700 62524 84756 62580
rect 84588 61292 84644 61348
rect 84588 60844 84644 60900
rect 85148 63922 85204 63924
rect 85148 63870 85150 63922
rect 85150 63870 85202 63922
rect 85202 63870 85204 63922
rect 85148 63868 85204 63870
rect 85484 64428 85540 64484
rect 85260 63084 85316 63140
rect 85372 63756 85428 63812
rect 85148 62636 85204 62692
rect 84028 60284 84084 60340
rect 83916 60172 83972 60228
rect 83804 57708 83860 57764
rect 82684 56700 82740 56756
rect 82572 55356 82628 55412
rect 82796 56588 82852 56644
rect 82908 57260 82964 57316
rect 82796 56082 82852 56084
rect 82796 56030 82798 56082
rect 82798 56030 82850 56082
rect 82850 56030 82852 56082
rect 82796 56028 82852 56030
rect 82572 54626 82628 54628
rect 82572 54574 82574 54626
rect 82574 54574 82626 54626
rect 82626 54574 82628 54626
rect 82572 54572 82628 54574
rect 82684 52332 82740 52388
rect 81228 51490 81284 51492
rect 81228 51438 81230 51490
rect 81230 51438 81282 51490
rect 81282 51438 81284 51490
rect 81228 51436 81284 51438
rect 81452 51490 81508 51492
rect 81452 51438 81454 51490
rect 81454 51438 81506 51490
rect 81506 51438 81508 51490
rect 81452 51436 81508 51438
rect 81900 51436 81956 51492
rect 81564 51100 81620 51156
rect 81564 50316 81620 50372
rect 81676 50428 81732 50484
rect 80556 50092 80612 50148
rect 81276 50202 81332 50204
rect 81276 50150 81278 50202
rect 81278 50150 81330 50202
rect 81330 50150 81332 50202
rect 81276 50148 81332 50150
rect 81380 50202 81436 50204
rect 81380 50150 81382 50202
rect 81382 50150 81434 50202
rect 81434 50150 81436 50202
rect 81380 50148 81436 50150
rect 81484 50202 81540 50204
rect 81484 50150 81486 50202
rect 81486 50150 81538 50202
rect 81538 50150 81540 50202
rect 81484 50148 81540 50150
rect 80444 49698 80500 49700
rect 80444 49646 80446 49698
rect 80446 49646 80498 49698
rect 80498 49646 80500 49698
rect 80444 49644 80500 49646
rect 80556 49532 80612 49588
rect 80108 48412 80164 48468
rect 81676 48972 81732 49028
rect 77756 42700 77812 42756
rect 77980 42700 78036 42756
rect 78540 42642 78596 42644
rect 78540 42590 78542 42642
rect 78542 42590 78594 42642
rect 78594 42590 78596 42642
rect 78540 42588 78596 42590
rect 77756 42028 77812 42084
rect 77420 41804 77476 41860
rect 78204 41858 78260 41860
rect 78204 41806 78206 41858
rect 78206 41806 78258 41858
rect 78258 41806 78260 41858
rect 78204 41804 78260 41806
rect 76524 41244 76580 41300
rect 76300 40962 76356 40964
rect 76300 40910 76302 40962
rect 76302 40910 76354 40962
rect 76354 40910 76356 40962
rect 76300 40908 76356 40910
rect 76412 39618 76468 39620
rect 76412 39566 76414 39618
rect 76414 39566 76466 39618
rect 76466 39566 76468 39618
rect 76412 39564 76468 39566
rect 76188 38946 76244 38948
rect 76188 38894 76190 38946
rect 76190 38894 76242 38946
rect 76242 38894 76244 38946
rect 76188 38892 76244 38894
rect 76524 37996 76580 38052
rect 76076 36540 76132 36596
rect 76412 36876 76468 36932
rect 74956 36204 75012 36260
rect 74732 35868 74788 35924
rect 76412 36204 76468 36260
rect 75292 35868 75348 35924
rect 76524 35810 76580 35812
rect 76524 35758 76526 35810
rect 76526 35758 76578 35810
rect 76578 35758 76580 35810
rect 76524 35756 76580 35758
rect 75516 34972 75572 35028
rect 76524 35026 76580 35028
rect 76524 34974 76526 35026
rect 76526 34974 76578 35026
rect 76578 34974 76580 35026
rect 76524 34972 76580 34974
rect 73724 33292 73780 33348
rect 74732 33346 74788 33348
rect 74732 33294 74734 33346
rect 74734 33294 74786 33346
rect 74786 33294 74788 33346
rect 74732 33292 74788 33294
rect 74284 33180 74340 33236
rect 73836 33068 73892 33124
rect 73836 32786 73892 32788
rect 73836 32734 73838 32786
rect 73838 32734 73890 32786
rect 73890 32734 73892 32786
rect 73836 32732 73892 32734
rect 74284 32786 74340 32788
rect 74284 32734 74286 32786
rect 74286 32734 74338 32786
rect 74338 32734 74340 32786
rect 74284 32732 74340 32734
rect 75516 32786 75572 32788
rect 75516 32734 75518 32786
rect 75518 32734 75570 32786
rect 75570 32734 75572 32786
rect 75516 32732 75572 32734
rect 76300 33346 76356 33348
rect 76300 33294 76302 33346
rect 76302 33294 76354 33346
rect 76354 33294 76356 33346
rect 76300 33292 76356 33294
rect 76188 32674 76244 32676
rect 76188 32622 76190 32674
rect 76190 32622 76242 32674
rect 76242 32622 76244 32674
rect 76188 32620 76244 32622
rect 76748 32786 76804 32788
rect 76748 32734 76750 32786
rect 76750 32734 76802 32786
rect 76802 32734 76804 32786
rect 76748 32732 76804 32734
rect 77308 41692 77364 41748
rect 77308 41074 77364 41076
rect 77308 41022 77310 41074
rect 77310 41022 77362 41074
rect 77362 41022 77364 41074
rect 77308 41020 77364 41022
rect 77196 40348 77252 40404
rect 77084 37884 77140 37940
rect 77308 39564 77364 39620
rect 77532 38780 77588 38836
rect 77756 40460 77812 40516
rect 78204 40460 78260 40516
rect 78316 38722 78372 38724
rect 78316 38670 78318 38722
rect 78318 38670 78370 38722
rect 78370 38670 78372 38722
rect 78316 38668 78372 38670
rect 79324 38722 79380 38724
rect 79324 38670 79326 38722
rect 79326 38670 79378 38722
rect 79378 38670 79380 38722
rect 79324 38668 79380 38670
rect 77756 38108 77812 38164
rect 77196 36876 77252 36932
rect 77532 36876 77588 36932
rect 77420 36540 77476 36596
rect 77084 34972 77140 35028
rect 77308 34914 77364 34916
rect 77308 34862 77310 34914
rect 77310 34862 77362 34914
rect 77362 34862 77364 34914
rect 77308 34860 77364 34862
rect 77308 32732 77364 32788
rect 77644 36594 77700 36596
rect 77644 36542 77646 36594
rect 77646 36542 77698 36594
rect 77698 36542 77700 36594
rect 77644 36540 77700 36542
rect 78988 38162 79044 38164
rect 78988 38110 78990 38162
rect 78990 38110 79042 38162
rect 79042 38110 79044 38162
rect 78988 38108 79044 38110
rect 77868 38050 77924 38052
rect 77868 37998 77870 38050
rect 77870 37998 77922 38050
rect 77922 37998 77924 38050
rect 77868 37996 77924 37998
rect 78540 38050 78596 38052
rect 78540 37998 78542 38050
rect 78542 37998 78594 38050
rect 78594 37998 78596 38050
rect 78540 37996 78596 37998
rect 77868 37378 77924 37380
rect 77868 37326 77870 37378
rect 77870 37326 77922 37378
rect 77922 37326 77924 37378
rect 77868 37324 77924 37326
rect 77756 34860 77812 34916
rect 77532 34300 77588 34356
rect 78764 34130 78820 34132
rect 78764 34078 78766 34130
rect 78766 34078 78818 34130
rect 78818 34078 78820 34130
rect 78764 34076 78820 34078
rect 77532 33292 77588 33348
rect 77868 33516 77924 33572
rect 81004 47570 81060 47572
rect 81004 47518 81006 47570
rect 81006 47518 81058 47570
rect 81058 47518 81060 47570
rect 81004 47516 81060 47518
rect 81004 46508 81060 46564
rect 80668 45778 80724 45780
rect 80668 45726 80670 45778
rect 80670 45726 80722 45778
rect 80722 45726 80724 45778
rect 80668 45724 80724 45726
rect 80668 45052 80724 45108
rect 80444 44156 80500 44212
rect 79548 42588 79604 42644
rect 80556 42812 80612 42868
rect 80556 41244 80612 41300
rect 80444 40402 80500 40404
rect 80444 40350 80446 40402
rect 80446 40350 80498 40402
rect 80498 40350 80500 40402
rect 80444 40348 80500 40350
rect 80108 38946 80164 38948
rect 80108 38894 80110 38946
rect 80110 38894 80162 38946
rect 80162 38894 80164 38946
rect 80108 38892 80164 38894
rect 79996 37996 80052 38052
rect 79996 37772 80052 37828
rect 79884 34242 79940 34244
rect 79884 34190 79886 34242
rect 79886 34190 79938 34242
rect 79938 34190 79940 34242
rect 79884 34188 79940 34190
rect 79436 33628 79492 33684
rect 80668 33292 80724 33348
rect 78988 32732 79044 32788
rect 77868 32674 77924 32676
rect 77868 32622 77870 32674
rect 77870 32622 77922 32674
rect 77922 32622 77924 32674
rect 77868 32620 77924 32622
rect 81276 48634 81332 48636
rect 81276 48582 81278 48634
rect 81278 48582 81330 48634
rect 81330 48582 81332 48634
rect 81276 48580 81332 48582
rect 81380 48634 81436 48636
rect 81380 48582 81382 48634
rect 81382 48582 81434 48634
rect 81434 48582 81436 48634
rect 81380 48580 81436 48582
rect 81484 48634 81540 48636
rect 81484 48582 81486 48634
rect 81486 48582 81538 48634
rect 81538 48582 81540 48634
rect 81484 48580 81540 48582
rect 82236 51436 82292 51492
rect 82012 51100 82068 51156
rect 82348 50092 82404 50148
rect 82236 49810 82292 49812
rect 82236 49758 82238 49810
rect 82238 49758 82290 49810
rect 82290 49758 82292 49810
rect 82236 49756 82292 49758
rect 81788 47628 81844 47684
rect 81676 47516 81732 47572
rect 82348 48354 82404 48356
rect 82348 48302 82350 48354
rect 82350 48302 82402 48354
rect 82402 48302 82404 48354
rect 82348 48300 82404 48302
rect 82236 47570 82292 47572
rect 82236 47518 82238 47570
rect 82238 47518 82290 47570
rect 82290 47518 82292 47570
rect 82236 47516 82292 47518
rect 81276 47066 81332 47068
rect 81276 47014 81278 47066
rect 81278 47014 81330 47066
rect 81330 47014 81332 47066
rect 81276 47012 81332 47014
rect 81380 47066 81436 47068
rect 81380 47014 81382 47066
rect 81382 47014 81434 47066
rect 81434 47014 81436 47066
rect 81380 47012 81436 47014
rect 81484 47066 81540 47068
rect 81484 47014 81486 47066
rect 81486 47014 81538 47066
rect 81538 47014 81540 47066
rect 81484 47012 81540 47014
rect 82572 46844 82628 46900
rect 81676 46562 81732 46564
rect 81676 46510 81678 46562
rect 81678 46510 81730 46562
rect 81730 46510 81732 46562
rect 81676 46508 81732 46510
rect 82236 46508 82292 46564
rect 82572 45890 82628 45892
rect 82572 45838 82574 45890
rect 82574 45838 82626 45890
rect 82626 45838 82628 45890
rect 82572 45836 82628 45838
rect 82796 50540 82852 50596
rect 82796 48300 82852 48356
rect 82796 45778 82852 45780
rect 82796 45726 82798 45778
rect 82798 45726 82850 45778
rect 82850 45726 82852 45778
rect 82796 45724 82852 45726
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 81116 45052 81172 45108
rect 81340 45106 81396 45108
rect 81340 45054 81342 45106
rect 81342 45054 81394 45106
rect 81394 45054 81396 45106
rect 81340 45052 81396 45054
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 81564 41074 81620 41076
rect 81564 41022 81566 41074
rect 81566 41022 81618 41074
rect 81618 41022 81620 41074
rect 81564 41020 81620 41022
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 81228 40402 81284 40404
rect 81228 40350 81230 40402
rect 81230 40350 81282 40402
rect 81282 40350 81284 40402
rect 81228 40348 81284 40350
rect 81340 39730 81396 39732
rect 81340 39678 81342 39730
rect 81342 39678 81394 39730
rect 81394 39678 81396 39730
rect 81340 39676 81396 39678
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 81452 39004 81508 39060
rect 81116 38892 81172 38948
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 81228 35922 81284 35924
rect 81228 35870 81230 35922
rect 81230 35870 81282 35922
rect 81282 35870 81284 35922
rect 81228 35868 81284 35870
rect 81788 41020 81844 41076
rect 82684 41074 82740 41076
rect 82684 41022 82686 41074
rect 82686 41022 82738 41074
rect 82738 41022 82740 41074
rect 82684 41020 82740 41022
rect 82460 40236 82516 40292
rect 82684 40124 82740 40180
rect 83468 57372 83524 57428
rect 83020 56588 83076 56644
rect 83244 55692 83300 55748
rect 83356 55356 83412 55412
rect 83020 54796 83076 54852
rect 83132 55244 83188 55300
rect 83020 53618 83076 53620
rect 83020 53566 83022 53618
rect 83022 53566 83074 53618
rect 83074 53566 83076 53618
rect 83020 53564 83076 53566
rect 83356 53788 83412 53844
rect 84028 58604 84084 58660
rect 84364 59948 84420 60004
rect 84476 59890 84532 59892
rect 84476 59838 84478 59890
rect 84478 59838 84530 59890
rect 84530 59838 84532 59890
rect 84476 59836 84532 59838
rect 84476 59052 84532 59108
rect 85484 61628 85540 61684
rect 85260 61570 85316 61572
rect 85260 61518 85262 61570
rect 85262 61518 85314 61570
rect 85314 61518 85316 61570
rect 85260 61516 85316 61518
rect 86268 70028 86324 70084
rect 86380 69804 86436 69860
rect 85708 69692 85764 69748
rect 86044 69522 86100 69524
rect 86044 69470 86046 69522
rect 86046 69470 86098 69522
rect 86098 69470 86100 69522
rect 86044 69468 86100 69470
rect 85820 68796 85876 68852
rect 86044 67730 86100 67732
rect 86044 67678 86046 67730
rect 86046 67678 86098 67730
rect 86098 67678 86100 67730
rect 86044 67676 86100 67678
rect 85820 67340 85876 67396
rect 86492 67282 86548 67284
rect 86492 67230 86494 67282
rect 86494 67230 86546 67282
rect 86546 67230 86548 67282
rect 86492 67228 86548 67230
rect 86492 66050 86548 66052
rect 86492 65998 86494 66050
rect 86494 65998 86546 66050
rect 86546 65998 86548 66050
rect 86492 65996 86548 65998
rect 86156 65660 86212 65716
rect 86716 67170 86772 67172
rect 86716 67118 86718 67170
rect 86718 67118 86770 67170
rect 86770 67118 86772 67170
rect 86716 67116 86772 67118
rect 86940 75628 86996 75684
rect 87052 75516 87108 75572
rect 87164 72546 87220 72548
rect 87164 72494 87166 72546
rect 87166 72494 87218 72546
rect 87218 72494 87220 72546
rect 87164 72492 87220 72494
rect 87164 70194 87220 70196
rect 87164 70142 87166 70194
rect 87166 70142 87218 70194
rect 87218 70142 87220 70194
rect 87164 70140 87220 70142
rect 87052 70028 87108 70084
rect 87164 69804 87220 69860
rect 86716 65602 86772 65604
rect 86716 65550 86718 65602
rect 86718 65550 86770 65602
rect 86770 65550 86772 65602
rect 86716 65548 86772 65550
rect 87052 66220 87108 66276
rect 86716 65266 86772 65268
rect 86716 65214 86718 65266
rect 86718 65214 86770 65266
rect 86770 65214 86772 65266
rect 86716 65212 86772 65214
rect 85932 63868 85988 63924
rect 85820 62860 85876 62916
rect 86044 63756 86100 63812
rect 86268 64092 86324 64148
rect 86268 63922 86324 63924
rect 86268 63870 86270 63922
rect 86270 63870 86322 63922
rect 86322 63870 86324 63922
rect 86268 63868 86324 63870
rect 86156 63250 86212 63252
rect 86156 63198 86158 63250
rect 86158 63198 86210 63250
rect 86210 63198 86212 63250
rect 86156 63196 86212 63198
rect 86268 63138 86324 63140
rect 86268 63086 86270 63138
rect 86270 63086 86322 63138
rect 86322 63086 86324 63138
rect 86268 63084 86324 63086
rect 86044 63026 86100 63028
rect 86044 62974 86046 63026
rect 86046 62974 86098 63026
rect 86098 62974 86100 63026
rect 86044 62972 86100 62974
rect 86044 62354 86100 62356
rect 86044 62302 86046 62354
rect 86046 62302 86098 62354
rect 86098 62302 86100 62354
rect 86044 62300 86100 62302
rect 86604 64092 86660 64148
rect 86604 62972 86660 63028
rect 86492 62354 86548 62356
rect 86492 62302 86494 62354
rect 86494 62302 86546 62354
rect 86546 62302 86548 62354
rect 86492 62300 86548 62302
rect 85708 62188 85764 62244
rect 86268 61740 86324 61796
rect 87388 68626 87444 68628
rect 87388 68574 87390 68626
rect 87390 68574 87442 68626
rect 87442 68574 87444 68626
rect 87388 68572 87444 68574
rect 87836 74114 87892 74116
rect 87836 74062 87838 74114
rect 87838 74062 87890 74114
rect 87890 74062 87892 74114
rect 87836 74060 87892 74062
rect 89292 86268 89348 86324
rect 88844 85314 88900 85316
rect 88844 85262 88846 85314
rect 88846 85262 88898 85314
rect 88898 85262 88900 85314
rect 88844 85260 88900 85262
rect 88172 85202 88228 85204
rect 88172 85150 88174 85202
rect 88174 85150 88226 85202
rect 88226 85150 88228 85202
rect 88172 85148 88228 85150
rect 89180 85202 89236 85204
rect 89180 85150 89182 85202
rect 89182 85150 89234 85202
rect 89234 85150 89236 85202
rect 89180 85148 89236 85150
rect 89292 84418 89348 84420
rect 89292 84366 89294 84418
rect 89294 84366 89346 84418
rect 89346 84366 89348 84418
rect 89292 84364 89348 84366
rect 88508 84306 88564 84308
rect 88508 84254 88510 84306
rect 88510 84254 88562 84306
rect 88562 84254 88564 84306
rect 88508 84252 88564 84254
rect 88284 84028 88340 84084
rect 88396 83468 88452 83524
rect 89404 84140 89460 84196
rect 88620 83746 88676 83748
rect 88620 83694 88622 83746
rect 88622 83694 88674 83746
rect 88674 83694 88676 83746
rect 88620 83692 88676 83694
rect 89516 84028 89572 84084
rect 88844 83244 88900 83300
rect 90188 84306 90244 84308
rect 90188 84254 90190 84306
rect 90190 84254 90242 84306
rect 90242 84254 90244 84306
rect 90188 84252 90244 84254
rect 89628 83244 89684 83300
rect 90524 84530 90580 84532
rect 90524 84478 90526 84530
rect 90526 84478 90578 84530
rect 90578 84478 90580 84530
rect 90524 84476 90580 84478
rect 92652 87388 92708 87444
rect 91532 86268 91588 86324
rect 91196 85036 91252 85092
rect 90748 83468 90804 83524
rect 91532 84194 91588 84196
rect 91532 84142 91534 84194
rect 91534 84142 91586 84194
rect 91586 84142 91588 84194
rect 91532 84140 91588 84142
rect 91532 83522 91588 83524
rect 91532 83470 91534 83522
rect 91534 83470 91586 83522
rect 91586 83470 91588 83522
rect 91532 83468 91588 83470
rect 92204 84476 92260 84532
rect 92204 83522 92260 83524
rect 92204 83470 92206 83522
rect 92206 83470 92258 83522
rect 92258 83470 92260 83522
rect 92204 83468 92260 83470
rect 92316 84978 92372 84980
rect 92316 84926 92318 84978
rect 92318 84926 92370 84978
rect 92370 84926 92372 84978
rect 92316 84924 92372 84926
rect 90412 82572 90468 82628
rect 90972 80668 91028 80724
rect 91196 80668 91252 80724
rect 88396 79884 88452 79940
rect 89628 79884 89684 79940
rect 89180 79826 89236 79828
rect 89180 79774 89182 79826
rect 89182 79774 89234 79826
rect 89234 79774 89236 79826
rect 89180 79772 89236 79774
rect 88396 78540 88452 78596
rect 90412 78764 90468 78820
rect 89516 78594 89572 78596
rect 89516 78542 89518 78594
rect 89518 78542 89570 78594
rect 89570 78542 89572 78594
rect 89516 78540 89572 78542
rect 89180 78034 89236 78036
rect 89180 77982 89182 78034
rect 89182 77982 89234 78034
rect 89234 77982 89236 78034
rect 89180 77980 89236 77982
rect 89516 78146 89572 78148
rect 89516 78094 89518 78146
rect 89518 78094 89570 78146
rect 89570 78094 89572 78146
rect 89516 78092 89572 78094
rect 89404 77308 89460 77364
rect 88284 74898 88340 74900
rect 88284 74846 88286 74898
rect 88286 74846 88338 74898
rect 88338 74846 88340 74898
rect 88284 74844 88340 74846
rect 89404 74898 89460 74900
rect 89404 74846 89406 74898
rect 89406 74846 89458 74898
rect 89458 74846 89460 74898
rect 89404 74844 89460 74846
rect 89068 74620 89124 74676
rect 91420 79660 91476 79716
rect 91868 79436 91924 79492
rect 91644 79324 91700 79380
rect 93548 85148 93604 85204
rect 93436 85090 93492 85092
rect 93436 85038 93438 85090
rect 93438 85038 93490 85090
rect 93490 85038 93492 85090
rect 93436 85036 93492 85038
rect 96636 88618 96692 88620
rect 96636 88566 96638 88618
rect 96638 88566 96690 88618
rect 96690 88566 96692 88618
rect 96636 88564 96692 88566
rect 96740 88618 96796 88620
rect 96740 88566 96742 88618
rect 96742 88566 96794 88618
rect 96794 88566 96796 88618
rect 96740 88564 96796 88566
rect 96844 88618 96900 88620
rect 96844 88566 96846 88618
rect 96846 88566 96898 88618
rect 96898 88566 96900 88618
rect 96844 88564 96900 88566
rect 94556 87442 94612 87444
rect 94556 87390 94558 87442
rect 94558 87390 94610 87442
rect 94610 87390 94612 87442
rect 94556 87388 94612 87390
rect 95116 87442 95172 87444
rect 95116 87390 95118 87442
rect 95118 87390 95170 87442
rect 95170 87390 95172 87442
rect 95116 87388 95172 87390
rect 96636 87050 96692 87052
rect 96636 86998 96638 87050
rect 96638 86998 96690 87050
rect 96690 86998 96692 87050
rect 96636 86996 96692 86998
rect 96740 87050 96796 87052
rect 96740 86998 96742 87050
rect 96742 86998 96794 87050
rect 96794 86998 96796 87050
rect 96740 86996 96796 86998
rect 96844 87050 96900 87052
rect 96844 86998 96846 87050
rect 96846 86998 96898 87050
rect 96898 86998 96900 87050
rect 96844 86996 96900 86998
rect 93772 84924 93828 84980
rect 94892 85148 94948 85204
rect 94444 84476 94500 84532
rect 92428 81730 92484 81732
rect 92428 81678 92430 81730
rect 92430 81678 92482 81730
rect 92482 81678 92484 81730
rect 92428 81676 92484 81678
rect 92204 81228 92260 81284
rect 92428 80668 92484 80724
rect 92540 79490 92596 79492
rect 92540 79438 92542 79490
rect 92542 79438 92594 79490
rect 92594 79438 92596 79490
rect 92540 79436 92596 79438
rect 94108 82012 94164 82068
rect 94220 84140 94276 84196
rect 93212 81058 93268 81060
rect 93212 81006 93214 81058
rect 93214 81006 93266 81058
rect 93266 81006 93268 81058
rect 93212 81004 93268 81006
rect 93100 80668 93156 80724
rect 93548 80668 93604 80724
rect 93324 80332 93380 80388
rect 94332 83634 94388 83636
rect 94332 83582 94334 83634
rect 94334 83582 94386 83634
rect 94386 83582 94388 83634
rect 94332 83580 94388 83582
rect 93884 81676 93940 81732
rect 94668 81058 94724 81060
rect 94668 81006 94670 81058
rect 94670 81006 94722 81058
rect 94722 81006 94724 81058
rect 94668 81004 94724 81006
rect 93884 80668 93940 80724
rect 94556 80668 94612 80724
rect 94332 80274 94388 80276
rect 94332 80222 94334 80274
rect 94334 80222 94386 80274
rect 94386 80222 94388 80274
rect 94332 80220 94388 80222
rect 93772 79660 93828 79716
rect 93996 79378 94052 79380
rect 93996 79326 93998 79378
rect 93998 79326 94050 79378
rect 94050 79326 94052 79378
rect 93996 79324 94052 79326
rect 90636 75180 90692 75236
rect 91420 75180 91476 75236
rect 89740 74786 89796 74788
rect 89740 74734 89742 74786
rect 89742 74734 89794 74786
rect 89794 74734 89796 74786
rect 89740 74732 89796 74734
rect 89516 74060 89572 74116
rect 89964 74620 90020 74676
rect 89964 74172 90020 74228
rect 89740 73948 89796 74004
rect 88060 70924 88116 70980
rect 88172 69244 88228 69300
rect 87724 68796 87780 68852
rect 88508 73330 88564 73332
rect 88508 73278 88510 73330
rect 88510 73278 88562 73330
rect 88562 73278 88564 73330
rect 88508 73276 88564 73278
rect 89404 73330 89460 73332
rect 89404 73278 89406 73330
rect 89406 73278 89458 73330
rect 89458 73278 89460 73330
rect 89404 73276 89460 73278
rect 90860 74732 90916 74788
rect 89180 71708 89236 71764
rect 89292 71148 89348 71204
rect 89404 70924 89460 70980
rect 89852 71762 89908 71764
rect 89852 71710 89854 71762
rect 89854 71710 89906 71762
rect 89906 71710 89908 71762
rect 89852 71708 89908 71710
rect 91756 74674 91812 74676
rect 91756 74622 91758 74674
rect 91758 74622 91810 74674
rect 91810 74622 91812 74674
rect 91756 74620 91812 74622
rect 91084 74172 91140 74228
rect 91308 74002 91364 74004
rect 91308 73950 91310 74002
rect 91310 73950 91362 74002
rect 91362 73950 91364 74002
rect 91308 73948 91364 73950
rect 90860 71148 90916 71204
rect 90860 70924 90916 70980
rect 89068 69410 89124 69412
rect 89068 69358 89070 69410
rect 89070 69358 89122 69410
rect 89122 69358 89124 69410
rect 89068 69356 89124 69358
rect 88844 69298 88900 69300
rect 88844 69246 88846 69298
rect 88846 69246 88898 69298
rect 88898 69246 88900 69298
rect 88844 69244 88900 69246
rect 88732 68796 88788 68852
rect 88508 68572 88564 68628
rect 89628 70194 89684 70196
rect 89628 70142 89630 70194
rect 89630 70142 89682 70194
rect 89682 70142 89684 70194
rect 89628 70140 89684 70142
rect 89628 69916 89684 69972
rect 89516 68684 89572 68740
rect 87500 67564 87556 67620
rect 88172 67228 88228 67284
rect 87724 67170 87780 67172
rect 87724 67118 87726 67170
rect 87726 67118 87778 67170
rect 87778 67118 87780 67170
rect 87724 67116 87780 67118
rect 88732 67116 88788 67172
rect 87836 67058 87892 67060
rect 87836 67006 87838 67058
rect 87838 67006 87890 67058
rect 87890 67006 87892 67058
rect 87836 67004 87892 67006
rect 87388 66274 87444 66276
rect 87388 66222 87390 66274
rect 87390 66222 87442 66274
rect 87442 66222 87444 66274
rect 87388 66220 87444 66222
rect 87948 66220 88004 66276
rect 87164 65996 87220 66052
rect 87612 63980 87668 64036
rect 87388 63868 87444 63924
rect 87052 63644 87108 63700
rect 86940 62748 86996 62804
rect 85820 61068 85876 61124
rect 84812 59948 84868 60004
rect 84812 58604 84868 58660
rect 85148 60060 85204 60116
rect 85260 59106 85316 59108
rect 85260 59054 85262 59106
rect 85262 59054 85314 59106
rect 85314 59054 85316 59106
rect 85260 59052 85316 59054
rect 84924 58268 84980 58324
rect 84476 57932 84532 57988
rect 83916 57260 83972 57316
rect 83804 57148 83860 57204
rect 83804 55020 83860 55076
rect 84028 55244 84084 55300
rect 84140 54572 84196 54628
rect 83916 54348 83972 54404
rect 84364 55020 84420 55076
rect 83580 53564 83636 53620
rect 83244 52332 83300 52388
rect 83804 50594 83860 50596
rect 83804 50542 83806 50594
rect 83806 50542 83858 50594
rect 83858 50542 83860 50594
rect 83804 50540 83860 50542
rect 84476 54572 84532 54628
rect 83580 49644 83636 49700
rect 83804 49756 83860 49812
rect 83020 49532 83076 49588
rect 84364 49810 84420 49812
rect 84364 49758 84366 49810
rect 84366 49758 84418 49810
rect 84418 49758 84420 49810
rect 84364 49756 84420 49758
rect 84140 49532 84196 49588
rect 83916 49420 83972 49476
rect 83804 48914 83860 48916
rect 83804 48862 83806 48914
rect 83806 48862 83858 48914
rect 83858 48862 83860 48914
rect 83804 48860 83860 48862
rect 83020 48802 83076 48804
rect 83020 48750 83022 48802
rect 83022 48750 83074 48802
rect 83074 48750 83076 48802
rect 83020 48748 83076 48750
rect 84364 49420 84420 49476
rect 84364 48972 84420 49028
rect 84700 57762 84756 57764
rect 84700 57710 84702 57762
rect 84702 57710 84754 57762
rect 84754 57710 84756 57762
rect 84700 57708 84756 57710
rect 85372 58492 85428 58548
rect 85596 60508 85652 60564
rect 85708 60732 85764 60788
rect 85596 60002 85652 60004
rect 85596 59950 85598 60002
rect 85598 59950 85650 60002
rect 85650 59950 85652 60002
rect 85596 59948 85652 59950
rect 86044 60002 86100 60004
rect 86044 59950 86046 60002
rect 86046 59950 86098 60002
rect 86098 59950 86100 60002
rect 86044 59948 86100 59950
rect 86828 62524 86884 62580
rect 87276 62636 87332 62692
rect 88060 65714 88116 65716
rect 88060 65662 88062 65714
rect 88062 65662 88114 65714
rect 88114 65662 88116 65714
rect 88060 65660 88116 65662
rect 88284 65548 88340 65604
rect 88956 67900 89012 67956
rect 88172 65490 88228 65492
rect 88172 65438 88174 65490
rect 88174 65438 88226 65490
rect 88226 65438 88228 65490
rect 88172 65436 88228 65438
rect 88844 65772 88900 65828
rect 88508 64988 88564 65044
rect 88396 64540 88452 64596
rect 88396 63308 88452 63364
rect 88396 63138 88452 63140
rect 88396 63086 88398 63138
rect 88398 63086 88450 63138
rect 88450 63086 88452 63138
rect 88396 63084 88452 63086
rect 87948 62636 88004 62692
rect 88060 62860 88116 62916
rect 87836 62466 87892 62468
rect 87836 62414 87838 62466
rect 87838 62414 87890 62466
rect 87890 62414 87892 62466
rect 87836 62412 87892 62414
rect 87612 61682 87668 61684
rect 87612 61630 87614 61682
rect 87614 61630 87666 61682
rect 87666 61630 87668 61682
rect 87612 61628 87668 61630
rect 87164 61346 87220 61348
rect 87164 61294 87166 61346
rect 87166 61294 87218 61346
rect 87218 61294 87220 61346
rect 87164 61292 87220 61294
rect 87052 60786 87108 60788
rect 87052 60734 87054 60786
rect 87054 60734 87106 60786
rect 87106 60734 87108 60786
rect 87052 60732 87108 60734
rect 86604 60620 86660 60676
rect 85148 55244 85204 55300
rect 85260 54626 85316 54628
rect 85260 54574 85262 54626
rect 85262 54574 85314 54626
rect 85314 54574 85316 54626
rect 85260 54572 85316 54574
rect 84700 54402 84756 54404
rect 84700 54350 84702 54402
rect 84702 54350 84754 54402
rect 84754 54350 84756 54402
rect 84700 54348 84756 54350
rect 85148 53618 85204 53620
rect 85148 53566 85150 53618
rect 85150 53566 85202 53618
rect 85202 53566 85204 53618
rect 85148 53564 85204 53566
rect 85260 52834 85316 52836
rect 85260 52782 85262 52834
rect 85262 52782 85314 52834
rect 85314 52782 85316 52834
rect 85260 52780 85316 52782
rect 84924 51212 84980 51268
rect 84588 50092 84644 50148
rect 84812 50540 84868 50596
rect 84812 49980 84868 50036
rect 84588 48860 84644 48916
rect 83132 46844 83188 46900
rect 84252 45836 84308 45892
rect 83356 45612 83412 45668
rect 83244 41074 83300 41076
rect 83244 41022 83246 41074
rect 83246 41022 83298 41074
rect 83298 41022 83300 41074
rect 83244 41020 83300 41022
rect 82908 39676 82964 39732
rect 82348 39618 82404 39620
rect 82348 39566 82350 39618
rect 82350 39566 82402 39618
rect 82402 39566 82404 39618
rect 82348 39564 82404 39566
rect 83244 39618 83300 39620
rect 83244 39566 83246 39618
rect 83246 39566 83298 39618
rect 83298 39566 83300 39618
rect 83244 39564 83300 39566
rect 82460 38780 82516 38836
rect 82236 37266 82292 37268
rect 82236 37214 82238 37266
rect 82238 37214 82290 37266
rect 82290 37214 82292 37266
rect 82236 37212 82292 37214
rect 81788 36764 81844 36820
rect 82572 39004 82628 39060
rect 83244 38108 83300 38164
rect 82908 37266 82964 37268
rect 82908 37214 82910 37266
rect 82910 37214 82962 37266
rect 82962 37214 82964 37266
rect 82908 37212 82964 37214
rect 83916 42028 83972 42084
rect 83804 40236 83860 40292
rect 83916 40402 83972 40404
rect 83916 40350 83918 40402
rect 83918 40350 83970 40402
rect 83970 40350 83972 40402
rect 83916 40348 83972 40350
rect 84140 42588 84196 42644
rect 83804 39676 83860 39732
rect 84476 47570 84532 47572
rect 84476 47518 84478 47570
rect 84478 47518 84530 47570
rect 84530 47518 84532 47570
rect 84476 47516 84532 47518
rect 84476 45778 84532 45780
rect 84476 45726 84478 45778
rect 84478 45726 84530 45778
rect 84530 45726 84532 45778
rect 84476 45724 84532 45726
rect 85260 50482 85316 50484
rect 85260 50430 85262 50482
rect 85262 50430 85314 50482
rect 85314 50430 85316 50482
rect 85260 50428 85316 50430
rect 85596 55132 85652 55188
rect 85484 52162 85540 52164
rect 85484 52110 85486 52162
rect 85486 52110 85538 52162
rect 85538 52110 85540 52162
rect 85484 52108 85540 52110
rect 85708 51884 85764 51940
rect 85036 49756 85092 49812
rect 85260 49644 85316 49700
rect 85036 48860 85092 48916
rect 85148 47628 85204 47684
rect 84924 45612 84980 45668
rect 84700 42028 84756 42084
rect 85596 49644 85652 49700
rect 86380 59052 86436 59108
rect 86492 58156 86548 58212
rect 85932 57650 85988 57652
rect 85932 57598 85934 57650
rect 85934 57598 85986 57650
rect 85986 57598 85988 57650
rect 85932 57596 85988 57598
rect 85932 55244 85988 55300
rect 86044 55186 86100 55188
rect 86044 55134 86046 55186
rect 86046 55134 86098 55186
rect 86098 55134 86100 55186
rect 86044 55132 86100 55134
rect 86380 53618 86436 53620
rect 86380 53566 86382 53618
rect 86382 53566 86434 53618
rect 86434 53566 86436 53618
rect 86380 53564 86436 53566
rect 86044 53452 86100 53508
rect 86044 52780 86100 52836
rect 86380 51884 86436 51940
rect 85820 50316 85876 50372
rect 85820 49420 85876 49476
rect 86828 57372 86884 57428
rect 86940 57260 86996 57316
rect 86604 56252 86660 56308
rect 85596 49026 85652 49028
rect 85596 48974 85598 49026
rect 85598 48974 85650 49026
rect 85650 48974 85652 49026
rect 85596 48972 85652 48974
rect 85708 48914 85764 48916
rect 85708 48862 85710 48914
rect 85710 48862 85762 48914
rect 85762 48862 85764 48914
rect 85708 48860 85764 48862
rect 85932 49026 85988 49028
rect 85932 48974 85934 49026
rect 85934 48974 85986 49026
rect 85986 48974 85988 49026
rect 85932 48972 85988 48974
rect 85820 47628 85876 47684
rect 85484 47404 85540 47460
rect 86492 49922 86548 49924
rect 86492 49870 86494 49922
rect 86494 49870 86546 49922
rect 86546 49870 86548 49922
rect 86492 49868 86548 49870
rect 86380 48972 86436 49028
rect 86268 48860 86324 48916
rect 86492 48076 86548 48132
rect 86044 47180 86100 47236
rect 85596 46732 85652 46788
rect 86268 46732 86324 46788
rect 85708 45890 85764 45892
rect 85708 45838 85710 45890
rect 85710 45838 85762 45890
rect 85762 45838 85764 45890
rect 85708 45836 85764 45838
rect 85932 45778 85988 45780
rect 85932 45726 85934 45778
rect 85934 45726 85986 45778
rect 85986 45726 85988 45778
rect 85932 45724 85988 45726
rect 86268 45778 86324 45780
rect 86268 45726 86270 45778
rect 86270 45726 86322 45778
rect 86322 45726 86324 45778
rect 86268 45724 86324 45726
rect 84252 41020 84308 41076
rect 84924 40236 84980 40292
rect 84140 40124 84196 40180
rect 86156 42754 86212 42756
rect 86156 42702 86158 42754
rect 86158 42702 86210 42754
rect 86210 42702 86212 42754
rect 86156 42700 86212 42702
rect 85260 42642 85316 42644
rect 85260 42590 85262 42642
rect 85262 42590 85314 42642
rect 85314 42590 85316 42642
rect 85260 42588 85316 42590
rect 86380 42642 86436 42644
rect 86380 42590 86382 42642
rect 86382 42590 86434 42642
rect 86434 42590 86436 42642
rect 86380 42588 86436 42590
rect 86828 54514 86884 54516
rect 86828 54462 86830 54514
rect 86830 54462 86882 54514
rect 86882 54462 86884 54514
rect 86828 54460 86884 54462
rect 86940 53618 86996 53620
rect 86940 53566 86942 53618
rect 86942 53566 86994 53618
rect 86994 53566 86996 53618
rect 86940 53564 86996 53566
rect 87052 53506 87108 53508
rect 87052 53454 87054 53506
rect 87054 53454 87106 53506
rect 87106 53454 87108 53506
rect 87052 53452 87108 53454
rect 87948 60508 88004 60564
rect 88172 62636 88228 62692
rect 87500 59388 87556 59444
rect 87276 58210 87332 58212
rect 87276 58158 87278 58210
rect 87278 58158 87330 58210
rect 87330 58158 87332 58210
rect 87276 58156 87332 58158
rect 87500 57596 87556 57652
rect 87388 57148 87444 57204
rect 87500 56082 87556 56084
rect 87500 56030 87502 56082
rect 87502 56030 87554 56082
rect 87554 56030 87556 56082
rect 87500 56028 87556 56030
rect 87500 54738 87556 54740
rect 87500 54686 87502 54738
rect 87502 54686 87554 54738
rect 87554 54686 87556 54738
rect 87500 54684 87556 54686
rect 87500 52162 87556 52164
rect 87500 52110 87502 52162
rect 87502 52110 87554 52162
rect 87554 52110 87556 52162
rect 87500 52108 87556 52110
rect 86940 51884 86996 51940
rect 87276 50316 87332 50372
rect 87836 58322 87892 58324
rect 87836 58270 87838 58322
rect 87838 58270 87890 58322
rect 87890 58270 87892 58322
rect 87836 58268 87892 58270
rect 88284 61516 88340 61572
rect 88620 64316 88676 64372
rect 88732 63196 88788 63252
rect 89068 67116 89124 67172
rect 89068 65772 89124 65828
rect 88956 65548 89012 65604
rect 89180 65490 89236 65492
rect 89180 65438 89182 65490
rect 89182 65438 89234 65490
rect 89234 65438 89236 65490
rect 89180 65436 89236 65438
rect 89516 65602 89572 65604
rect 89516 65550 89518 65602
rect 89518 65550 89570 65602
rect 89570 65550 89572 65602
rect 89516 65548 89572 65550
rect 89404 64764 89460 64820
rect 88956 63308 89012 63364
rect 88620 62300 88676 62356
rect 89068 62412 89124 62468
rect 89292 63922 89348 63924
rect 89292 63870 89294 63922
rect 89294 63870 89346 63922
rect 89346 63870 89348 63922
rect 89292 63868 89348 63870
rect 89516 63644 89572 63700
rect 89516 63308 89572 63364
rect 89628 63084 89684 63140
rect 89292 62466 89348 62468
rect 89292 62414 89294 62466
rect 89294 62414 89346 62466
rect 89346 62414 89348 62466
rect 89292 62412 89348 62414
rect 89516 62300 89572 62356
rect 88508 60620 88564 60676
rect 89628 61570 89684 61572
rect 89628 61518 89630 61570
rect 89630 61518 89682 61570
rect 89682 61518 89684 61570
rect 89628 61516 89684 61518
rect 91308 71036 91364 71092
rect 90300 69356 90356 69412
rect 90524 68908 90580 68964
rect 90188 68684 90244 68740
rect 90188 68348 90244 68404
rect 90972 69916 91028 69972
rect 91196 68626 91252 68628
rect 91196 68574 91198 68626
rect 91198 68574 91250 68626
rect 91250 68574 91252 68626
rect 91196 68572 91252 68574
rect 90972 68012 91028 68068
rect 90860 67004 90916 67060
rect 91644 74226 91700 74228
rect 91644 74174 91646 74226
rect 91646 74174 91698 74226
rect 91698 74174 91700 74226
rect 91644 74172 91700 74174
rect 91756 73330 91812 73332
rect 91756 73278 91758 73330
rect 91758 73278 91810 73330
rect 91810 73278 91812 73330
rect 91756 73276 91812 73278
rect 91756 72380 91812 72436
rect 91644 69298 91700 69300
rect 91644 69246 91646 69298
rect 91646 69246 91698 69298
rect 91698 69246 91700 69298
rect 91644 69244 91700 69246
rect 90972 66332 91028 66388
rect 90972 66162 91028 66164
rect 90972 66110 90974 66162
rect 90974 66110 91026 66162
rect 91026 66110 91028 66162
rect 90972 66108 91028 66110
rect 90076 65996 90132 66052
rect 90860 66050 90916 66052
rect 90860 65998 90862 66050
rect 90862 65998 90914 66050
rect 90914 65998 90916 66050
rect 90860 65996 90916 65998
rect 90188 65772 90244 65828
rect 90860 65714 90916 65716
rect 90860 65662 90862 65714
rect 90862 65662 90914 65714
rect 90914 65662 90916 65714
rect 90860 65660 90916 65662
rect 90300 65602 90356 65604
rect 90300 65550 90302 65602
rect 90302 65550 90354 65602
rect 90354 65550 90356 65602
rect 90300 65548 90356 65550
rect 90636 65548 90692 65604
rect 90188 64764 90244 64820
rect 90076 63196 90132 63252
rect 90300 64146 90356 64148
rect 90300 64094 90302 64146
rect 90302 64094 90354 64146
rect 90354 64094 90356 64146
rect 90300 64092 90356 64094
rect 90412 63868 90468 63924
rect 90300 62972 90356 63028
rect 89740 60786 89796 60788
rect 89740 60734 89742 60786
rect 89742 60734 89794 60786
rect 89794 60734 89796 60786
rect 89740 60732 89796 60734
rect 89292 60508 89348 60564
rect 89068 59948 89124 60004
rect 88396 59724 88452 59780
rect 88844 59724 88900 59780
rect 88172 59276 88228 59332
rect 88508 58546 88564 58548
rect 88508 58494 88510 58546
rect 88510 58494 88562 58546
rect 88562 58494 88564 58546
rect 88508 58492 88564 58494
rect 87724 57260 87780 57316
rect 88172 57372 88228 57428
rect 87948 57260 88004 57316
rect 86940 49532 86996 49588
rect 87276 49756 87332 49812
rect 87500 49810 87556 49812
rect 87500 49758 87502 49810
rect 87502 49758 87554 49810
rect 87554 49758 87556 49810
rect 87500 49756 87556 49758
rect 88620 57650 88676 57652
rect 88620 57598 88622 57650
rect 88622 57598 88674 57650
rect 88674 57598 88676 57650
rect 88620 57596 88676 57598
rect 88508 57260 88564 57316
rect 88620 57148 88676 57204
rect 88620 56306 88676 56308
rect 88620 56254 88622 56306
rect 88622 56254 88674 56306
rect 88674 56254 88676 56306
rect 88620 56252 88676 56254
rect 88284 56194 88340 56196
rect 88284 56142 88286 56194
rect 88286 56142 88338 56194
rect 88338 56142 88340 56194
rect 88284 56140 88340 56142
rect 87836 54572 87892 54628
rect 88172 54514 88228 54516
rect 88172 54462 88174 54514
rect 88174 54462 88226 54514
rect 88226 54462 88228 54514
rect 88172 54460 88228 54462
rect 88284 54236 88340 54292
rect 87836 49810 87892 49812
rect 87836 49758 87838 49810
rect 87838 49758 87890 49810
rect 87890 49758 87892 49810
rect 87836 49756 87892 49758
rect 87724 47964 87780 48020
rect 87836 49532 87892 49588
rect 87724 47458 87780 47460
rect 87724 47406 87726 47458
rect 87726 47406 87778 47458
rect 87778 47406 87780 47458
rect 87724 47404 87780 47406
rect 87612 47234 87668 47236
rect 87612 47182 87614 47234
rect 87614 47182 87666 47234
rect 87666 47182 87668 47234
rect 87612 47180 87668 47182
rect 88284 49980 88340 50036
rect 88284 49810 88340 49812
rect 88284 49758 88286 49810
rect 88286 49758 88338 49810
rect 88338 49758 88340 49810
rect 88284 49756 88340 49758
rect 88396 49586 88452 49588
rect 88396 49534 88398 49586
rect 88398 49534 88450 49586
rect 88450 49534 88452 49586
rect 88396 49532 88452 49534
rect 88060 47964 88116 48020
rect 87724 45724 87780 45780
rect 86604 42476 86660 42532
rect 86716 42700 86772 42756
rect 85820 40236 85876 40292
rect 83580 38108 83636 38164
rect 84476 39004 84532 39060
rect 84252 38162 84308 38164
rect 84252 38110 84254 38162
rect 84254 38110 84306 38162
rect 84306 38110 84308 38162
rect 84252 38108 84308 38110
rect 83804 37100 83860 37156
rect 81788 35868 81844 35924
rect 81788 35308 81844 35364
rect 81676 34748 81732 34804
rect 82124 34860 82180 34916
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 81116 33628 81172 33684
rect 82348 34188 82404 34244
rect 82124 33628 82180 33684
rect 82460 34076 82516 34132
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 81340 32786 81396 32788
rect 81340 32734 81342 32786
rect 81342 32734 81394 32786
rect 81394 32734 81396 32786
rect 81340 32732 81396 32734
rect 76972 25228 77028 25284
rect 73388 12684 73444 12740
rect 69132 3330 69188 3332
rect 69132 3278 69134 3330
rect 69134 3278 69186 3330
rect 69186 3278 69188 3330
rect 69132 3276 69188 3278
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 81276 25114 81332 25116
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 82348 30940 82404 30996
rect 85148 39004 85204 39060
rect 87948 39730 88004 39732
rect 87948 39678 87950 39730
rect 87950 39678 88002 39730
rect 88002 39678 88004 39730
rect 87948 39676 88004 39678
rect 85820 39058 85876 39060
rect 85820 39006 85822 39058
rect 85822 39006 85874 39058
rect 85874 39006 85876 39058
rect 85820 39004 85876 39006
rect 84588 37154 84644 37156
rect 84588 37102 84590 37154
rect 84590 37102 84642 37154
rect 84642 37102 84644 37154
rect 84588 37100 84644 37102
rect 86716 36540 86772 36596
rect 82908 35196 82964 35252
rect 82684 34914 82740 34916
rect 82684 34862 82686 34914
rect 82686 34862 82738 34914
rect 82738 34862 82740 34914
rect 82684 34860 82740 34862
rect 83244 34802 83300 34804
rect 83244 34750 83246 34802
rect 83246 34750 83298 34802
rect 83298 34750 83300 34802
rect 83244 34748 83300 34750
rect 82796 33346 82852 33348
rect 82796 33294 82798 33346
rect 82798 33294 82850 33346
rect 82850 33294 82852 33346
rect 82796 33292 82852 33294
rect 84924 36428 84980 36484
rect 84924 35756 84980 35812
rect 86156 35810 86212 35812
rect 86156 35758 86158 35810
rect 86158 35758 86210 35810
rect 86210 35758 86212 35810
rect 86156 35756 86212 35758
rect 87052 36594 87108 36596
rect 87052 36542 87054 36594
rect 87054 36542 87106 36594
rect 87106 36542 87108 36594
rect 87052 36540 87108 36542
rect 84252 34914 84308 34916
rect 84252 34862 84254 34914
rect 84254 34862 84306 34914
rect 84306 34862 84308 34914
rect 84252 34860 84308 34862
rect 85596 34860 85652 34916
rect 84476 34802 84532 34804
rect 84476 34750 84478 34802
rect 84478 34750 84530 34802
rect 84530 34750 84532 34802
rect 84476 34748 84532 34750
rect 85148 34412 85204 34468
rect 83916 33852 83972 33908
rect 82908 32732 82964 32788
rect 83692 32732 83748 32788
rect 83132 30994 83188 30996
rect 83132 30942 83134 30994
rect 83134 30942 83186 30994
rect 83186 30942 83188 30994
rect 83132 30940 83188 30942
rect 84364 32732 84420 32788
rect 86044 34802 86100 34804
rect 86044 34750 86046 34802
rect 86046 34750 86098 34802
rect 86098 34750 86100 34802
rect 86044 34748 86100 34750
rect 85932 34412 85988 34468
rect 87500 34412 87556 34468
rect 86492 34188 86548 34244
rect 85820 34076 85876 34132
rect 86604 34130 86660 34132
rect 86604 34078 86606 34130
rect 86606 34078 86658 34130
rect 86658 34078 86660 34130
rect 86604 34076 86660 34078
rect 86940 34076 86996 34132
rect 86716 33628 86772 33684
rect 85596 33180 85652 33236
rect 86044 32786 86100 32788
rect 86044 32734 86046 32786
rect 86046 32734 86098 32786
rect 86098 32734 86100 32786
rect 86044 32732 86100 32734
rect 85596 32620 85652 32676
rect 84588 30828 84644 30884
rect 83692 29484 83748 29540
rect 83244 29426 83300 29428
rect 83244 29374 83246 29426
rect 83246 29374 83298 29426
rect 83298 29374 83300 29426
rect 83244 29372 83300 29374
rect 85148 29538 85204 29540
rect 85148 29486 85150 29538
rect 85150 29486 85202 29538
rect 85202 29486 85204 29538
rect 85148 29484 85204 29486
rect 87948 35756 88004 35812
rect 87612 34188 87668 34244
rect 87276 33906 87332 33908
rect 87276 33854 87278 33906
rect 87278 33854 87330 33906
rect 87330 33854 87332 33906
rect 87276 33852 87332 33854
rect 88172 47628 88228 47684
rect 88620 48130 88676 48132
rect 88620 48078 88622 48130
rect 88622 48078 88674 48130
rect 88674 48078 88676 48130
rect 88620 48076 88676 48078
rect 88508 47180 88564 47236
rect 88620 45948 88676 46004
rect 88284 42530 88340 42532
rect 88284 42478 88286 42530
rect 88286 42478 88338 42530
rect 88338 42478 88340 42530
rect 88284 42476 88340 42478
rect 88732 42140 88788 42196
rect 88172 40236 88228 40292
rect 88508 42028 88564 42084
rect 89404 59778 89460 59780
rect 89404 59726 89406 59778
rect 89406 59726 89458 59778
rect 89458 59726 89460 59778
rect 89404 59724 89460 59726
rect 89292 58268 89348 58324
rect 89516 57148 89572 57204
rect 89852 59388 89908 59444
rect 89628 56364 89684 56420
rect 89292 54738 89348 54740
rect 89292 54686 89294 54738
rect 89294 54686 89346 54738
rect 89346 54686 89348 54738
rect 89292 54684 89348 54686
rect 89628 55692 89684 55748
rect 89516 54626 89572 54628
rect 89516 54574 89518 54626
rect 89518 54574 89570 54626
rect 89570 54574 89572 54626
rect 89516 54572 89572 54574
rect 89852 54684 89908 54740
rect 89404 53788 89460 53844
rect 89516 54124 89572 54180
rect 90076 58492 90132 58548
rect 90188 58940 90244 58996
rect 90076 56252 90132 56308
rect 90076 54124 90132 54180
rect 89964 54012 90020 54068
rect 90300 56194 90356 56196
rect 90300 56142 90302 56194
rect 90302 56142 90354 56194
rect 90354 56142 90356 56194
rect 90300 56140 90356 56142
rect 91980 74284 92036 74340
rect 92316 75010 92372 75012
rect 92316 74958 92318 75010
rect 92318 74958 92370 75010
rect 92370 74958 92372 75010
rect 92316 74956 92372 74958
rect 92092 74732 92148 74788
rect 92428 74620 92484 74676
rect 93548 75740 93604 75796
rect 93212 74956 93268 75012
rect 94332 78876 94388 78932
rect 94444 77980 94500 78036
rect 94444 76972 94500 77028
rect 93772 74732 93828 74788
rect 93548 74620 93604 74676
rect 92540 74172 92596 74228
rect 91868 71596 91924 71652
rect 91980 71148 92036 71204
rect 92316 73276 92372 73332
rect 93100 74284 93156 74340
rect 93660 73442 93716 73444
rect 93660 73390 93662 73442
rect 93662 73390 93714 73442
rect 93714 73390 93716 73442
rect 93660 73388 93716 73390
rect 92540 72268 92596 72324
rect 91980 70978 92036 70980
rect 91980 70926 91982 70978
rect 91982 70926 92034 70978
rect 92034 70926 92036 70978
rect 91980 70924 92036 70926
rect 92988 71148 93044 71204
rect 93660 71090 93716 71092
rect 93660 71038 93662 71090
rect 93662 71038 93714 71090
rect 93714 71038 93716 71090
rect 93660 71036 93716 71038
rect 93100 70978 93156 70980
rect 93100 70926 93102 70978
rect 93102 70926 93154 70978
rect 93154 70926 93156 70978
rect 93100 70924 93156 70926
rect 93212 69298 93268 69300
rect 93212 69246 93214 69298
rect 93214 69246 93266 69298
rect 93266 69246 93268 69298
rect 93212 69244 93268 69246
rect 93436 68908 93492 68964
rect 91532 66220 91588 66276
rect 91868 68572 91924 68628
rect 91420 66162 91476 66164
rect 91420 66110 91422 66162
rect 91422 66110 91474 66162
rect 91474 66110 91476 66162
rect 91420 66108 91476 66110
rect 91308 65996 91364 66052
rect 90748 64818 90804 64820
rect 90748 64766 90750 64818
rect 90750 64766 90802 64818
rect 90802 64766 90804 64818
rect 90748 64764 90804 64766
rect 90748 63644 90804 63700
rect 90860 63756 90916 63812
rect 90636 58546 90692 58548
rect 90636 58494 90638 58546
rect 90638 58494 90690 58546
rect 90690 58494 90692 58546
rect 90636 58492 90692 58494
rect 90524 56306 90580 56308
rect 90524 56254 90526 56306
rect 90526 56254 90578 56306
rect 90578 56254 90580 56306
rect 90524 56252 90580 56254
rect 90636 55692 90692 55748
rect 91308 64092 91364 64148
rect 91196 63644 91252 63700
rect 91196 63138 91252 63140
rect 91196 63086 91198 63138
rect 91198 63086 91250 63138
rect 91250 63086 91252 63138
rect 91196 63084 91252 63086
rect 91532 62188 91588 62244
rect 92092 68348 92148 68404
rect 93548 67954 93604 67956
rect 93548 67902 93550 67954
rect 93550 67902 93602 67954
rect 93602 67902 93604 67954
rect 93548 67900 93604 67902
rect 91868 67004 91924 67060
rect 91868 65548 91924 65604
rect 92204 63250 92260 63252
rect 92204 63198 92206 63250
rect 92206 63198 92258 63250
rect 92258 63198 92260 63250
rect 92204 63196 92260 63198
rect 91756 62914 91812 62916
rect 91756 62862 91758 62914
rect 91758 62862 91810 62914
rect 91810 62862 91812 62914
rect 91756 62860 91812 62862
rect 92988 63922 93044 63924
rect 92988 63870 92990 63922
rect 92990 63870 93042 63922
rect 93042 63870 93044 63922
rect 92988 63868 93044 63870
rect 92540 63756 92596 63812
rect 92316 62860 92372 62916
rect 93100 62412 93156 62468
rect 92316 62354 92372 62356
rect 92316 62302 92318 62354
rect 92318 62302 92370 62354
rect 92370 62302 92372 62354
rect 92316 62300 92372 62302
rect 92540 61404 92596 61460
rect 91644 60956 91700 61012
rect 91868 61180 91924 61236
rect 91420 58434 91476 58436
rect 91420 58382 91422 58434
rect 91422 58382 91474 58434
rect 91474 58382 91476 58434
rect 91420 58380 91476 58382
rect 91756 58380 91812 58436
rect 92428 60844 92484 60900
rect 92204 60508 92260 60564
rect 91980 58380 92036 58436
rect 91420 57650 91476 57652
rect 91420 57598 91422 57650
rect 91422 57598 91474 57650
rect 91474 57598 91476 57650
rect 91420 57596 91476 57598
rect 90300 54626 90356 54628
rect 90300 54574 90302 54626
rect 90302 54574 90354 54626
rect 90354 54574 90356 54626
rect 90300 54572 90356 54574
rect 90412 54514 90468 54516
rect 90412 54462 90414 54514
rect 90414 54462 90466 54514
rect 90466 54462 90468 54514
rect 90412 54460 90468 54462
rect 90188 53004 90244 53060
rect 90300 54012 90356 54068
rect 90076 52946 90132 52948
rect 90076 52894 90078 52946
rect 90078 52894 90130 52946
rect 90130 52894 90132 52946
rect 90076 52892 90132 52894
rect 89628 51884 89684 51940
rect 89964 51266 90020 51268
rect 89964 51214 89966 51266
rect 89966 51214 90018 51266
rect 90018 51214 90020 51266
rect 89964 51212 90020 51214
rect 90188 51772 90244 51828
rect 88956 49756 89012 49812
rect 89068 50428 89124 50484
rect 89068 49084 89124 49140
rect 89068 46002 89124 46004
rect 89068 45950 89070 46002
rect 89070 45950 89122 46002
rect 89122 45950 89124 46002
rect 89068 45948 89124 45950
rect 88172 36540 88228 36596
rect 88060 34636 88116 34692
rect 87836 33628 87892 33684
rect 88508 37826 88564 37828
rect 88508 37774 88510 37826
rect 88510 37774 88562 37826
rect 88562 37774 88564 37826
rect 88508 37772 88564 37774
rect 88844 40572 88900 40628
rect 89292 50482 89348 50484
rect 89292 50430 89294 50482
rect 89294 50430 89346 50482
rect 89346 50430 89348 50482
rect 89292 50428 89348 50430
rect 90076 50652 90132 50708
rect 90076 50316 90132 50372
rect 90188 50428 90244 50484
rect 90300 49922 90356 49924
rect 90300 49870 90302 49922
rect 90302 49870 90354 49922
rect 90354 49870 90356 49922
rect 90300 49868 90356 49870
rect 89292 49810 89348 49812
rect 89292 49758 89294 49810
rect 89294 49758 89346 49810
rect 89346 49758 89348 49810
rect 89292 49756 89348 49758
rect 89292 48748 89348 48804
rect 89740 47180 89796 47236
rect 89740 45890 89796 45892
rect 89740 45838 89742 45890
rect 89742 45838 89794 45890
rect 89794 45838 89796 45890
rect 89740 45836 89796 45838
rect 89852 47068 89908 47124
rect 90860 54738 90916 54740
rect 90860 54686 90862 54738
rect 90862 54686 90914 54738
rect 90914 54686 90916 54738
rect 90860 54684 90916 54686
rect 91084 54626 91140 54628
rect 91084 54574 91086 54626
rect 91086 54574 91138 54626
rect 91138 54574 91140 54626
rect 91084 54572 91140 54574
rect 91196 54514 91252 54516
rect 91196 54462 91198 54514
rect 91198 54462 91250 54514
rect 91250 54462 91252 54514
rect 91196 54460 91252 54462
rect 90748 53788 90804 53844
rect 90860 53676 90916 53732
rect 91196 53788 91252 53844
rect 91644 54236 91700 54292
rect 91084 50594 91140 50596
rect 91084 50542 91086 50594
rect 91086 50542 91138 50594
rect 91138 50542 91140 50594
rect 91084 50540 91140 50542
rect 90748 49868 90804 49924
rect 91196 50316 91252 50372
rect 93212 62188 93268 62244
rect 93212 61682 93268 61684
rect 93212 61630 93214 61682
rect 93214 61630 93266 61682
rect 93266 61630 93268 61682
rect 93212 61628 93268 61630
rect 94332 75010 94388 75012
rect 94332 74958 94334 75010
rect 94334 74958 94386 75010
rect 94386 74958 94388 75010
rect 94332 74956 94388 74958
rect 93996 73948 94052 74004
rect 93996 73388 94052 73444
rect 94108 72322 94164 72324
rect 94108 72270 94110 72322
rect 94110 72270 94162 72322
rect 94162 72270 94164 72322
rect 94108 72268 94164 72270
rect 93996 67058 94052 67060
rect 93996 67006 93998 67058
rect 93998 67006 94050 67058
rect 94050 67006 94052 67058
rect 93996 67004 94052 67006
rect 93772 66892 93828 66948
rect 94108 66780 94164 66836
rect 94108 66386 94164 66388
rect 94108 66334 94110 66386
rect 94110 66334 94162 66386
rect 94162 66334 94164 66386
rect 94108 66332 94164 66334
rect 94332 65490 94388 65492
rect 94332 65438 94334 65490
rect 94334 65438 94386 65490
rect 94386 65438 94388 65490
rect 94332 65436 94388 65438
rect 93772 64988 93828 65044
rect 94220 64988 94276 65044
rect 93660 64482 93716 64484
rect 93660 64430 93662 64482
rect 93662 64430 93714 64482
rect 93714 64430 93716 64482
rect 93660 64428 93716 64430
rect 96636 85482 96692 85484
rect 96636 85430 96638 85482
rect 96638 85430 96690 85482
rect 96690 85430 96692 85482
rect 96636 85428 96692 85430
rect 96740 85482 96796 85484
rect 96740 85430 96742 85482
rect 96742 85430 96794 85482
rect 96794 85430 96796 85482
rect 96740 85428 96796 85430
rect 96844 85482 96900 85484
rect 96844 85430 96846 85482
rect 96846 85430 96898 85482
rect 96898 85430 96900 85482
rect 96844 85428 96900 85430
rect 95564 84476 95620 84532
rect 95788 83580 95844 83636
rect 96348 84418 96404 84420
rect 96348 84366 96350 84418
rect 96350 84366 96402 84418
rect 96402 84366 96404 84418
rect 96348 84364 96404 84366
rect 95788 82124 95844 82180
rect 94892 80386 94948 80388
rect 94892 80334 94894 80386
rect 94894 80334 94946 80386
rect 94946 80334 94948 80386
rect 94892 80332 94948 80334
rect 94892 79714 94948 79716
rect 94892 79662 94894 79714
rect 94894 79662 94946 79714
rect 94946 79662 94948 79714
rect 94892 79660 94948 79662
rect 96236 83468 96292 83524
rect 96636 83914 96692 83916
rect 96636 83862 96638 83914
rect 96638 83862 96690 83914
rect 96690 83862 96692 83914
rect 96636 83860 96692 83862
rect 96740 83914 96796 83916
rect 96740 83862 96742 83914
rect 96742 83862 96794 83914
rect 96794 83862 96796 83914
rect 96740 83860 96796 83862
rect 96844 83914 96900 83916
rect 96844 83862 96846 83914
rect 96846 83862 96898 83914
rect 96898 83862 96900 83914
rect 96844 83860 96900 83862
rect 96636 82346 96692 82348
rect 96636 82294 96638 82346
rect 96638 82294 96690 82346
rect 96690 82294 96692 82346
rect 96636 82292 96692 82294
rect 96740 82346 96796 82348
rect 96740 82294 96742 82346
rect 96742 82294 96794 82346
rect 96794 82294 96796 82346
rect 96740 82292 96796 82294
rect 96844 82346 96900 82348
rect 96844 82294 96846 82346
rect 96846 82294 96898 82346
rect 96898 82294 96900 82346
rect 96844 82292 96900 82294
rect 97356 82066 97412 82068
rect 97356 82014 97358 82066
rect 97358 82014 97410 82066
rect 97410 82014 97412 82066
rect 97356 82012 97412 82014
rect 95564 81058 95620 81060
rect 95564 81006 95566 81058
rect 95566 81006 95618 81058
rect 95618 81006 95620 81058
rect 95564 81004 95620 81006
rect 95340 80444 95396 80500
rect 95340 79884 95396 79940
rect 95452 80556 95508 80612
rect 95228 79660 95284 79716
rect 94780 76972 94836 77028
rect 97244 81058 97300 81060
rect 97244 81006 97246 81058
rect 97246 81006 97298 81058
rect 97298 81006 97300 81058
rect 97244 81004 97300 81006
rect 96636 80778 96692 80780
rect 96636 80726 96638 80778
rect 96638 80726 96690 80778
rect 96690 80726 96692 80778
rect 96636 80724 96692 80726
rect 96740 80778 96796 80780
rect 96740 80726 96742 80778
rect 96742 80726 96794 80778
rect 96794 80726 96796 80778
rect 96740 80724 96796 80726
rect 96844 80778 96900 80780
rect 96844 80726 96846 80778
rect 96846 80726 96898 80778
rect 96898 80726 96900 80778
rect 96844 80724 96900 80726
rect 96124 80556 96180 80612
rect 95788 80220 95844 80276
rect 95676 79772 95732 79828
rect 97244 79826 97300 79828
rect 97244 79774 97246 79826
rect 97246 79774 97298 79826
rect 97298 79774 97300 79826
rect 97244 79772 97300 79774
rect 96124 79714 96180 79716
rect 96124 79662 96126 79714
rect 96126 79662 96178 79714
rect 96178 79662 96180 79714
rect 96124 79660 96180 79662
rect 96348 79548 96404 79604
rect 95564 78540 95620 78596
rect 96636 79210 96692 79212
rect 96636 79158 96638 79210
rect 96638 79158 96690 79210
rect 96690 79158 96692 79210
rect 96636 79156 96692 79158
rect 96740 79210 96796 79212
rect 96740 79158 96742 79210
rect 96742 79158 96794 79210
rect 96794 79158 96796 79210
rect 96740 79156 96796 79158
rect 96844 79210 96900 79212
rect 96844 79158 96846 79210
rect 96846 79158 96898 79210
rect 96898 79158 96900 79210
rect 96844 79156 96900 79158
rect 95228 78034 95284 78036
rect 95228 77982 95230 78034
rect 95230 77982 95282 78034
rect 95282 77982 95284 78034
rect 95228 77980 95284 77982
rect 95004 77026 95060 77028
rect 95004 76974 95006 77026
rect 95006 76974 95058 77026
rect 95058 76974 95060 77026
rect 95004 76972 95060 76974
rect 96636 77642 96692 77644
rect 96636 77590 96638 77642
rect 96638 77590 96690 77642
rect 96690 77590 96692 77642
rect 96636 77588 96692 77590
rect 96740 77642 96796 77644
rect 96740 77590 96742 77642
rect 96742 77590 96794 77642
rect 96794 77590 96796 77642
rect 96740 77588 96796 77590
rect 96844 77642 96900 77644
rect 96844 77590 96846 77642
rect 96846 77590 96898 77642
rect 96898 77590 96900 77642
rect 96844 77588 96900 77590
rect 96012 76972 96068 77028
rect 97132 76972 97188 77028
rect 96636 76074 96692 76076
rect 96636 76022 96638 76074
rect 96638 76022 96690 76074
rect 96690 76022 96692 76074
rect 96636 76020 96692 76022
rect 96740 76074 96796 76076
rect 96740 76022 96742 76074
rect 96742 76022 96794 76074
rect 96794 76022 96796 76074
rect 96740 76020 96796 76022
rect 96844 76074 96900 76076
rect 96844 76022 96846 76074
rect 96846 76022 96898 76074
rect 96898 76022 96900 76074
rect 96844 76020 96900 76022
rect 95340 75794 95396 75796
rect 95340 75742 95342 75794
rect 95342 75742 95394 75794
rect 95394 75742 95396 75794
rect 95340 75740 95396 75742
rect 94892 75628 94948 75684
rect 94556 74956 94612 75012
rect 96012 75682 96068 75684
rect 96012 75630 96014 75682
rect 96014 75630 96066 75682
rect 96066 75630 96068 75682
rect 96012 75628 96068 75630
rect 96348 74786 96404 74788
rect 96348 74734 96350 74786
rect 96350 74734 96402 74786
rect 96402 74734 96404 74786
rect 96348 74732 96404 74734
rect 96636 74506 96692 74508
rect 96636 74454 96638 74506
rect 96638 74454 96690 74506
rect 96690 74454 96692 74506
rect 96636 74452 96692 74454
rect 96740 74506 96796 74508
rect 96740 74454 96742 74506
rect 96742 74454 96794 74506
rect 96794 74454 96796 74506
rect 96740 74452 96796 74454
rect 96844 74506 96900 74508
rect 96844 74454 96846 74506
rect 96846 74454 96898 74506
rect 96898 74454 96900 74506
rect 96844 74452 96900 74454
rect 96348 74172 96404 74228
rect 95788 73948 95844 74004
rect 97132 73948 97188 74004
rect 95228 73330 95284 73332
rect 95228 73278 95230 73330
rect 95230 73278 95282 73330
rect 95282 73278 95284 73330
rect 95228 73276 95284 73278
rect 94668 72492 94724 72548
rect 96636 72938 96692 72940
rect 96636 72886 96638 72938
rect 96638 72886 96690 72938
rect 96690 72886 96692 72938
rect 96636 72884 96692 72886
rect 96740 72938 96796 72940
rect 96740 72886 96742 72938
rect 96742 72886 96794 72938
rect 96794 72886 96796 72938
rect 96740 72884 96796 72886
rect 96844 72938 96900 72940
rect 96844 72886 96846 72938
rect 96846 72886 96898 72938
rect 96898 72886 96900 72938
rect 96844 72884 96900 72886
rect 94556 72380 94612 72436
rect 95564 71650 95620 71652
rect 95564 71598 95566 71650
rect 95566 71598 95618 71650
rect 95618 71598 95620 71650
rect 95564 71596 95620 71598
rect 96636 71370 96692 71372
rect 96636 71318 96638 71370
rect 96638 71318 96690 71370
rect 96690 71318 96692 71370
rect 96636 71316 96692 71318
rect 96740 71370 96796 71372
rect 96740 71318 96742 71370
rect 96742 71318 96794 71370
rect 96794 71318 96796 71370
rect 96740 71316 96796 71318
rect 96844 71370 96900 71372
rect 96844 71318 96846 71370
rect 96846 71318 96898 71370
rect 96898 71318 96900 71370
rect 96844 71316 96900 71318
rect 95004 71036 95060 71092
rect 96460 71090 96516 71092
rect 96460 71038 96462 71090
rect 96462 71038 96514 71090
rect 96514 71038 96516 71090
rect 96460 71036 96516 71038
rect 95452 70252 95508 70308
rect 94892 69522 94948 69524
rect 94892 69470 94894 69522
rect 94894 69470 94946 69522
rect 94946 69470 94948 69522
rect 94892 69468 94948 69470
rect 94668 67788 94724 67844
rect 95116 70082 95172 70084
rect 95116 70030 95118 70082
rect 95118 70030 95170 70082
rect 95170 70030 95172 70082
rect 95116 70028 95172 70030
rect 95116 67900 95172 67956
rect 95340 69468 95396 69524
rect 95676 70476 95732 70532
rect 95676 69468 95732 69524
rect 96012 69468 96068 69524
rect 96460 70194 96516 70196
rect 96460 70142 96462 70194
rect 96462 70142 96514 70194
rect 96514 70142 96516 70194
rect 96460 70140 96516 70142
rect 97132 70082 97188 70084
rect 97132 70030 97134 70082
rect 97134 70030 97186 70082
rect 97186 70030 97188 70082
rect 97132 70028 97188 70030
rect 96636 69802 96692 69804
rect 96636 69750 96638 69802
rect 96638 69750 96690 69802
rect 96690 69750 96692 69802
rect 96636 69748 96692 69750
rect 96740 69802 96796 69804
rect 96740 69750 96742 69802
rect 96742 69750 96794 69802
rect 96794 69750 96796 69802
rect 96740 69748 96796 69750
rect 96844 69802 96900 69804
rect 96844 69750 96846 69802
rect 96846 69750 96898 69802
rect 96898 69750 96900 69802
rect 96844 69748 96900 69750
rect 97020 69522 97076 69524
rect 97020 69470 97022 69522
rect 97022 69470 97074 69522
rect 97074 69470 97076 69522
rect 97020 69468 97076 69470
rect 96636 68234 96692 68236
rect 96636 68182 96638 68234
rect 96638 68182 96690 68234
rect 96690 68182 96692 68234
rect 96636 68180 96692 68182
rect 96740 68234 96796 68236
rect 96740 68182 96742 68234
rect 96742 68182 96794 68234
rect 96794 68182 96796 68234
rect 96740 68180 96796 68182
rect 96844 68234 96900 68236
rect 96844 68182 96846 68234
rect 96846 68182 96898 68234
rect 96898 68182 96900 68234
rect 96844 68180 96900 68182
rect 96348 67842 96404 67844
rect 96348 67790 96350 67842
rect 96350 67790 96402 67842
rect 96402 67790 96404 67842
rect 96348 67788 96404 67790
rect 97356 67842 97412 67844
rect 97356 67790 97358 67842
rect 97358 67790 97410 67842
rect 97410 67790 97412 67842
rect 97356 67788 97412 67790
rect 95452 67116 95508 67172
rect 96348 67170 96404 67172
rect 96348 67118 96350 67170
rect 96350 67118 96402 67170
rect 96402 67118 96404 67170
rect 96348 67116 96404 67118
rect 95228 66780 95284 66836
rect 95788 67004 95844 67060
rect 95340 65436 95396 65492
rect 94444 64428 94500 64484
rect 93436 64146 93492 64148
rect 93436 64094 93438 64146
rect 93438 64094 93490 64146
rect 93490 64094 93492 64146
rect 93436 64092 93492 64094
rect 94556 64146 94612 64148
rect 94556 64094 94558 64146
rect 94558 64094 94610 64146
rect 94610 64094 94612 64146
rect 94556 64092 94612 64094
rect 95004 63084 95060 63140
rect 93660 62636 93716 62692
rect 93324 61180 93380 61236
rect 94220 62914 94276 62916
rect 94220 62862 94222 62914
rect 94222 62862 94274 62914
rect 94274 62862 94276 62914
rect 94220 62860 94276 62862
rect 94332 62636 94388 62692
rect 94108 60508 94164 60564
rect 94332 60002 94388 60004
rect 94332 59950 94334 60002
rect 94334 59950 94386 60002
rect 94386 59950 94388 60002
rect 94332 59948 94388 59950
rect 94444 59330 94500 59332
rect 94444 59278 94446 59330
rect 94446 59278 94498 59330
rect 94498 59278 94500 59330
rect 94444 59276 94500 59278
rect 95116 62636 95172 62692
rect 95564 64988 95620 65044
rect 95452 61628 95508 61684
rect 95564 64428 95620 64484
rect 95676 62636 95732 62692
rect 94668 61458 94724 61460
rect 94668 61406 94670 61458
rect 94670 61406 94722 61458
rect 94722 61406 94724 61458
rect 94668 61404 94724 61406
rect 92316 57708 92372 57764
rect 92204 57650 92260 57652
rect 92204 57598 92206 57650
rect 92206 57598 92258 57650
rect 92258 57598 92260 57650
rect 92204 57596 92260 57598
rect 92428 57596 92484 57652
rect 91868 56588 91924 56644
rect 92204 56252 92260 56308
rect 91980 55916 92036 55972
rect 91756 51996 91812 52052
rect 91868 53900 91924 53956
rect 91532 50482 91588 50484
rect 91532 50430 91534 50482
rect 91534 50430 91586 50482
rect 91586 50430 91588 50482
rect 91532 50428 91588 50430
rect 92316 55916 92372 55972
rect 92316 55692 92372 55748
rect 92204 55244 92260 55300
rect 92092 54402 92148 54404
rect 92092 54350 92094 54402
rect 92094 54350 92146 54402
rect 92146 54350 92148 54402
rect 92092 54348 92148 54350
rect 92092 53900 92148 53956
rect 92204 53788 92260 53844
rect 92316 54796 92372 54852
rect 92540 53676 92596 53732
rect 94892 58322 94948 58324
rect 94892 58270 94894 58322
rect 94894 58270 94946 58322
rect 94946 58270 94948 58322
rect 94892 58268 94948 58270
rect 92764 57762 92820 57764
rect 92764 57710 92766 57762
rect 92766 57710 92818 57762
rect 92818 57710 92820 57762
rect 92764 57708 92820 57710
rect 92764 54796 92820 54852
rect 93100 56924 93156 56980
rect 94332 57762 94388 57764
rect 94332 57710 94334 57762
rect 94334 57710 94386 57762
rect 94386 57710 94388 57762
rect 94332 57708 94388 57710
rect 93324 56642 93380 56644
rect 93324 56590 93326 56642
rect 93326 56590 93378 56642
rect 93378 56590 93380 56642
rect 93324 56588 93380 56590
rect 93100 56364 93156 56420
rect 93660 57650 93716 57652
rect 93660 57598 93662 57650
rect 93662 57598 93714 57650
rect 93714 57598 93716 57650
rect 93660 57596 93716 57598
rect 93660 56812 93716 56868
rect 94332 56866 94388 56868
rect 94332 56814 94334 56866
rect 94334 56814 94386 56866
rect 94386 56814 94388 56866
rect 94332 56812 94388 56814
rect 93884 56588 93940 56644
rect 93436 55692 93492 55748
rect 93548 55804 93604 55860
rect 93548 55298 93604 55300
rect 93548 55246 93550 55298
rect 93550 55246 93602 55298
rect 93602 55246 93604 55298
rect 93548 55244 93604 55246
rect 93548 54796 93604 54852
rect 94332 55804 94388 55860
rect 95340 57708 95396 57764
rect 95004 56978 95060 56980
rect 95004 56926 95006 56978
rect 95006 56926 95058 56978
rect 95058 56926 95060 56978
rect 95004 56924 95060 56926
rect 96908 67004 96964 67060
rect 96012 66946 96068 66948
rect 96012 66894 96014 66946
rect 96014 66894 96066 66946
rect 96066 66894 96068 66946
rect 96012 66892 96068 66894
rect 97132 66946 97188 66948
rect 97132 66894 97134 66946
rect 97134 66894 97186 66946
rect 97186 66894 97188 66946
rect 97132 66892 97188 66894
rect 96124 66780 96180 66836
rect 96636 66666 96692 66668
rect 96636 66614 96638 66666
rect 96638 66614 96690 66666
rect 96690 66614 96692 66666
rect 96636 66612 96692 66614
rect 96740 66666 96796 66668
rect 96740 66614 96742 66666
rect 96742 66614 96794 66666
rect 96794 66614 96796 66666
rect 96740 66612 96796 66614
rect 96844 66666 96900 66668
rect 96844 66614 96846 66666
rect 96846 66614 96898 66666
rect 96898 66614 96900 66666
rect 96844 66612 96900 66614
rect 97804 84364 97860 84420
rect 97692 80444 97748 80500
rect 97804 80556 97860 80612
rect 97580 79602 97636 79604
rect 97580 79550 97582 79602
rect 97582 79550 97634 79602
rect 97634 79550 97636 79602
rect 97580 79548 97636 79550
rect 97804 78540 97860 78596
rect 97804 74226 97860 74228
rect 97804 74174 97806 74226
rect 97806 74174 97858 74226
rect 97858 74174 97860 74226
rect 97804 74172 97860 74174
rect 98252 75068 98308 75124
rect 97580 73330 97636 73332
rect 97580 73278 97582 73330
rect 97582 73278 97634 73330
rect 97634 73278 97636 73330
rect 97580 73276 97636 73278
rect 97692 72546 97748 72548
rect 97692 72494 97694 72546
rect 97694 72494 97746 72546
rect 97746 72494 97748 72546
rect 97692 72492 97748 72494
rect 97692 70140 97748 70196
rect 98028 67788 98084 67844
rect 97580 66780 97636 66836
rect 97468 66444 97524 66500
rect 96348 65602 96404 65604
rect 96348 65550 96350 65602
rect 96350 65550 96402 65602
rect 96402 65550 96404 65602
rect 96348 65548 96404 65550
rect 97580 65548 97636 65604
rect 96636 65098 96692 65100
rect 96636 65046 96638 65098
rect 96638 65046 96690 65098
rect 96690 65046 96692 65098
rect 96636 65044 96692 65046
rect 96740 65098 96796 65100
rect 96740 65046 96742 65098
rect 96742 65046 96794 65098
rect 96794 65046 96796 65098
rect 96740 65044 96796 65046
rect 96844 65098 96900 65100
rect 96844 65046 96846 65098
rect 96846 65046 96898 65098
rect 96898 65046 96900 65098
rect 96844 65044 96900 65046
rect 97132 64706 97188 64708
rect 97132 64654 97134 64706
rect 97134 64654 97186 64706
rect 97186 64654 97188 64706
rect 97132 64652 97188 64654
rect 97692 64652 97748 64708
rect 96348 64092 96404 64148
rect 96636 63530 96692 63532
rect 96636 63478 96638 63530
rect 96638 63478 96690 63530
rect 96690 63478 96692 63530
rect 96636 63476 96692 63478
rect 96740 63530 96796 63532
rect 96740 63478 96742 63530
rect 96742 63478 96794 63530
rect 96794 63478 96796 63530
rect 96740 63476 96796 63478
rect 96844 63530 96900 63532
rect 96844 63478 96846 63530
rect 96846 63478 96898 63530
rect 96898 63478 96900 63530
rect 96844 63476 96900 63478
rect 96460 63084 96516 63140
rect 96348 62300 96404 62356
rect 97020 62860 97076 62916
rect 96636 61962 96692 61964
rect 96636 61910 96638 61962
rect 96638 61910 96690 61962
rect 96690 61910 96692 61962
rect 96636 61908 96692 61910
rect 96740 61962 96796 61964
rect 96740 61910 96742 61962
rect 96742 61910 96794 61962
rect 96794 61910 96796 61962
rect 96740 61908 96796 61910
rect 96844 61962 96900 61964
rect 96844 61910 96846 61962
rect 96846 61910 96898 61962
rect 96898 61910 96900 61962
rect 96844 61908 96900 61910
rect 97244 62636 97300 62692
rect 96636 60394 96692 60396
rect 96636 60342 96638 60394
rect 96638 60342 96690 60394
rect 96690 60342 96692 60394
rect 96636 60340 96692 60342
rect 96740 60394 96796 60396
rect 96740 60342 96742 60394
rect 96742 60342 96794 60394
rect 96794 60342 96796 60394
rect 96740 60340 96796 60342
rect 96844 60394 96900 60396
rect 96844 60342 96846 60394
rect 96846 60342 96898 60394
rect 96898 60342 96900 60394
rect 96844 60340 96900 60342
rect 98140 60732 98196 60788
rect 97692 60002 97748 60004
rect 97692 59950 97694 60002
rect 97694 59950 97746 60002
rect 97746 59950 97748 60002
rect 97692 59948 97748 59950
rect 97356 59890 97412 59892
rect 97356 59838 97358 59890
rect 97358 59838 97410 59890
rect 97410 59838 97412 59890
rect 97356 59836 97412 59838
rect 98028 59890 98084 59892
rect 98028 59838 98030 59890
rect 98030 59838 98082 59890
rect 98082 59838 98084 59890
rect 98028 59836 98084 59838
rect 95564 59330 95620 59332
rect 95564 59278 95566 59330
rect 95566 59278 95618 59330
rect 95618 59278 95620 59330
rect 95564 59276 95620 59278
rect 96636 58826 96692 58828
rect 96636 58774 96638 58826
rect 96638 58774 96690 58826
rect 96690 58774 96692 58826
rect 96636 58772 96692 58774
rect 96740 58826 96796 58828
rect 96740 58774 96742 58826
rect 96742 58774 96794 58826
rect 96794 58774 96796 58826
rect 96740 58772 96796 58774
rect 96844 58826 96900 58828
rect 96844 58774 96846 58826
rect 96846 58774 96898 58826
rect 96898 58774 96900 58826
rect 96844 58772 96900 58774
rect 96124 57820 96180 57876
rect 97580 58268 97636 58324
rect 96460 58044 96516 58100
rect 96908 58044 96964 58100
rect 97356 58044 97412 58100
rect 96636 57258 96692 57260
rect 96636 57206 96638 57258
rect 96638 57206 96690 57258
rect 96690 57206 96692 57258
rect 96636 57204 96692 57206
rect 96740 57258 96796 57260
rect 96740 57206 96742 57258
rect 96742 57206 96794 57258
rect 96794 57206 96796 57258
rect 96740 57204 96796 57206
rect 96844 57258 96900 57260
rect 96844 57206 96846 57258
rect 96846 57206 96898 57258
rect 96898 57206 96900 57258
rect 96844 57204 96900 57206
rect 95564 56588 95620 56644
rect 96236 55804 96292 55860
rect 92876 53900 92932 53956
rect 93100 53900 93156 53956
rect 93660 54626 93716 54628
rect 93660 54574 93662 54626
rect 93662 54574 93714 54626
rect 93714 54574 93716 54626
rect 93660 54572 93716 54574
rect 93660 54012 93716 54068
rect 94444 54236 94500 54292
rect 95004 54236 95060 54292
rect 94780 53676 94836 53732
rect 94108 53564 94164 53620
rect 91868 50652 91924 50708
rect 91868 50482 91924 50484
rect 91868 50430 91870 50482
rect 91870 50430 91922 50482
rect 91922 50430 91924 50482
rect 91868 50428 91924 50430
rect 91196 49980 91252 50036
rect 90972 47516 91028 47572
rect 91420 46844 91476 46900
rect 89628 45612 89684 45668
rect 90076 44044 90132 44100
rect 89740 42754 89796 42756
rect 89740 42702 89742 42754
rect 89742 42702 89794 42754
rect 89794 42702 89796 42754
rect 89740 42700 89796 42702
rect 89292 42476 89348 42532
rect 89292 40626 89348 40628
rect 89292 40574 89294 40626
rect 89294 40574 89346 40626
rect 89346 40574 89348 40626
rect 89292 40572 89348 40574
rect 89740 41356 89796 41412
rect 89628 41186 89684 41188
rect 89628 41134 89630 41186
rect 89630 41134 89682 41186
rect 89682 41134 89684 41186
rect 89628 41132 89684 41134
rect 90860 45948 90916 46004
rect 90524 45890 90580 45892
rect 90524 45838 90526 45890
rect 90526 45838 90578 45890
rect 90578 45838 90580 45890
rect 90524 45836 90580 45838
rect 91308 46002 91364 46004
rect 91308 45950 91310 46002
rect 91310 45950 91362 46002
rect 91362 45950 91364 46002
rect 91308 45948 91364 45950
rect 91196 45836 91252 45892
rect 90748 45778 90804 45780
rect 90748 45726 90750 45778
rect 90750 45726 90802 45778
rect 90802 45726 90804 45778
rect 90748 45724 90804 45726
rect 90636 44098 90692 44100
rect 90636 44046 90638 44098
rect 90638 44046 90690 44098
rect 90690 44046 90692 44098
rect 90636 44044 90692 44046
rect 91308 44044 91364 44100
rect 90076 42812 90132 42868
rect 89964 42140 90020 42196
rect 89852 41244 89908 41300
rect 90300 41410 90356 41412
rect 90300 41358 90302 41410
rect 90302 41358 90354 41410
rect 90354 41358 90356 41410
rect 90300 41356 90356 41358
rect 90412 41244 90468 41300
rect 90188 38892 90244 38948
rect 89516 37996 89572 38052
rect 89404 37324 89460 37380
rect 89292 37154 89348 37156
rect 89292 37102 89294 37154
rect 89294 37102 89346 37154
rect 89346 37102 89348 37154
rect 89292 37100 89348 37102
rect 88732 36540 88788 36596
rect 88508 35810 88564 35812
rect 88508 35758 88510 35810
rect 88510 35758 88562 35810
rect 88562 35758 88564 35810
rect 88508 35756 88564 35758
rect 90300 37100 90356 37156
rect 89964 35810 90020 35812
rect 89964 35758 89966 35810
rect 89966 35758 90018 35810
rect 90018 35758 90020 35810
rect 89964 35756 90020 35758
rect 89516 34860 89572 34916
rect 88396 34076 88452 34132
rect 88620 34636 88676 34692
rect 88172 32732 88228 32788
rect 89180 34076 89236 34132
rect 89404 34130 89460 34132
rect 89404 34078 89406 34130
rect 89406 34078 89458 34130
rect 89458 34078 89460 34130
rect 89404 34076 89460 34078
rect 89516 33628 89572 33684
rect 87388 32674 87444 32676
rect 87388 32622 87390 32674
rect 87390 32622 87442 32674
rect 87442 32622 87444 32674
rect 87388 32620 87444 32622
rect 86044 30882 86100 30884
rect 86044 30830 86046 30882
rect 86046 30830 86098 30882
rect 86098 30830 86100 30882
rect 86044 30828 86100 30830
rect 89292 31890 89348 31892
rect 89292 31838 89294 31890
rect 89294 31838 89346 31890
rect 89346 31838 89348 31890
rect 89292 31836 89348 31838
rect 87052 30828 87108 30884
rect 85372 29426 85428 29428
rect 85372 29374 85374 29426
rect 85374 29374 85426 29426
rect 85426 29374 85428 29426
rect 85372 29372 85428 29374
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 77532 2828 77588 2884
rect 69020 2716 69076 2772
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 90748 41132 90804 41188
rect 91420 43484 91476 43540
rect 91308 41186 91364 41188
rect 91308 41134 91310 41186
rect 91310 41134 91362 41186
rect 91362 41134 91364 41186
rect 91308 41132 91364 41134
rect 90636 39676 90692 39732
rect 91756 49644 91812 49700
rect 92428 50594 92484 50596
rect 92428 50542 92430 50594
rect 92430 50542 92482 50594
rect 92482 50542 92484 50594
rect 92428 50540 92484 50542
rect 92540 50428 92596 50484
rect 92652 49756 92708 49812
rect 92204 48300 92260 48356
rect 92092 47570 92148 47572
rect 92092 47518 92094 47570
rect 92094 47518 92146 47570
rect 92146 47518 92148 47570
rect 92092 47516 92148 47518
rect 91980 46844 92036 46900
rect 92428 46002 92484 46004
rect 92428 45950 92430 46002
rect 92430 45950 92482 46002
rect 92482 45950 92484 46002
rect 92428 45948 92484 45950
rect 92540 45724 92596 45780
rect 91980 45666 92036 45668
rect 91980 45614 91982 45666
rect 91982 45614 92034 45666
rect 92034 45614 92036 45666
rect 91980 45612 92036 45614
rect 91980 44322 92036 44324
rect 91980 44270 91982 44322
rect 91982 44270 92034 44322
rect 92034 44270 92036 44322
rect 91980 44268 92036 44270
rect 93996 52892 94052 52948
rect 92988 50540 93044 50596
rect 92876 48354 92932 48356
rect 92876 48302 92878 48354
rect 92878 48302 92930 48354
rect 92930 48302 92932 48354
rect 92876 48300 92932 48302
rect 93212 51548 93268 51604
rect 93324 50370 93380 50372
rect 93324 50318 93326 50370
rect 93326 50318 93378 50370
rect 93378 50318 93380 50370
rect 93324 50316 93380 50318
rect 94668 53058 94724 53060
rect 94668 53006 94670 53058
rect 94670 53006 94722 53058
rect 94722 53006 94724 53058
rect 94668 53004 94724 53006
rect 94556 52946 94612 52948
rect 94556 52894 94558 52946
rect 94558 52894 94610 52946
rect 94610 52894 94612 52946
rect 94556 52892 94612 52894
rect 94332 52162 94388 52164
rect 94332 52110 94334 52162
rect 94334 52110 94386 52162
rect 94386 52110 94388 52162
rect 94332 52108 94388 52110
rect 93996 51548 94052 51604
rect 94108 51772 94164 51828
rect 93996 51100 94052 51156
rect 93884 50428 93940 50484
rect 93772 48914 93828 48916
rect 93772 48862 93774 48914
rect 93774 48862 93826 48914
rect 93826 48862 93828 48914
rect 93772 48860 93828 48862
rect 93660 48242 93716 48244
rect 93660 48190 93662 48242
rect 93662 48190 93714 48242
rect 93714 48190 93716 48242
rect 93660 48188 93716 48190
rect 93436 48076 93492 48132
rect 93212 47346 93268 47348
rect 93212 47294 93214 47346
rect 93214 47294 93266 47346
rect 93266 47294 93268 47346
rect 93212 47292 93268 47294
rect 93324 47180 93380 47236
rect 93548 47404 93604 47460
rect 93660 47292 93716 47348
rect 93100 46396 93156 46452
rect 94892 52668 94948 52724
rect 94668 51548 94724 51604
rect 95004 51436 95060 51492
rect 94108 50204 94164 50260
rect 94332 50370 94388 50372
rect 94332 50318 94334 50370
rect 94334 50318 94386 50370
rect 94386 50318 94388 50370
rect 94332 50316 94388 50318
rect 94892 50204 94948 50260
rect 94220 48188 94276 48244
rect 94332 48130 94388 48132
rect 94332 48078 94334 48130
rect 94334 48078 94386 48130
rect 94386 48078 94388 48130
rect 94332 48076 94388 48078
rect 94444 47964 94500 48020
rect 94108 47292 94164 47348
rect 93996 47068 94052 47124
rect 94220 47068 94276 47124
rect 93884 46956 93940 47012
rect 93772 46898 93828 46900
rect 93772 46846 93774 46898
rect 93774 46846 93826 46898
rect 93826 46846 93828 46898
rect 93772 46844 93828 46846
rect 93660 46508 93716 46564
rect 92988 45948 93044 46004
rect 93324 45836 93380 45892
rect 93100 45666 93156 45668
rect 93100 45614 93102 45666
rect 93102 45614 93154 45666
rect 93154 45614 93156 45666
rect 93100 45612 93156 45614
rect 92316 42700 92372 42756
rect 92652 43538 92708 43540
rect 92652 43486 92654 43538
rect 92654 43486 92706 43538
rect 92706 43486 92708 43538
rect 92652 43484 92708 43486
rect 92428 42530 92484 42532
rect 92428 42478 92430 42530
rect 92430 42478 92482 42530
rect 92482 42478 92484 42530
rect 92428 42476 92484 42478
rect 92652 42028 92708 42084
rect 92652 41804 92708 41860
rect 92428 41074 92484 41076
rect 92428 41022 92430 41074
rect 92430 41022 92482 41074
rect 92482 41022 92484 41074
rect 92428 41020 92484 41022
rect 91532 38892 91588 38948
rect 91196 38834 91252 38836
rect 91196 38782 91198 38834
rect 91198 38782 91250 38834
rect 91250 38782 91252 38834
rect 91196 38780 91252 38782
rect 89852 34300 89908 34356
rect 91644 38050 91700 38052
rect 91644 37998 91646 38050
rect 91646 37998 91698 38050
rect 91698 37998 91700 38050
rect 91644 37996 91700 37998
rect 90972 37772 91028 37828
rect 91420 37378 91476 37380
rect 91420 37326 91422 37378
rect 91422 37326 91474 37378
rect 91474 37326 91476 37378
rect 91420 37324 91476 37326
rect 91980 37324 92036 37380
rect 90972 36540 91028 36596
rect 91644 36988 91700 37044
rect 92764 36988 92820 37044
rect 91644 34914 91700 34916
rect 91644 34862 91646 34914
rect 91646 34862 91698 34914
rect 91698 34862 91700 34914
rect 91644 34860 91700 34862
rect 90972 34412 91028 34468
rect 91980 34188 92036 34244
rect 92988 42140 93044 42196
rect 94332 46956 94388 47012
rect 93212 42754 93268 42756
rect 93212 42702 93214 42754
rect 93214 42702 93266 42754
rect 93266 42702 93268 42754
rect 93212 42700 93268 42702
rect 93548 44322 93604 44324
rect 93548 44270 93550 44322
rect 93550 44270 93602 44322
rect 93602 44270 93604 44322
rect 93548 44268 93604 44270
rect 93548 41244 93604 41300
rect 93660 40460 93716 40516
rect 94892 49922 94948 49924
rect 94892 49870 94894 49922
rect 94894 49870 94946 49922
rect 94946 49870 94948 49922
rect 94892 49868 94948 49870
rect 94780 49644 94836 49700
rect 94780 48188 94836 48244
rect 97244 55970 97300 55972
rect 97244 55918 97246 55970
rect 97246 55918 97298 55970
rect 97298 55918 97300 55970
rect 97244 55916 97300 55918
rect 97020 55804 97076 55860
rect 96636 55690 96692 55692
rect 96636 55638 96638 55690
rect 96638 55638 96690 55690
rect 96690 55638 96692 55690
rect 96636 55636 96692 55638
rect 96740 55690 96796 55692
rect 96740 55638 96742 55690
rect 96742 55638 96794 55690
rect 96794 55638 96796 55690
rect 96740 55636 96796 55638
rect 96844 55690 96900 55692
rect 96844 55638 96846 55690
rect 96846 55638 96898 55690
rect 96898 55638 96900 55690
rect 96844 55636 96900 55638
rect 97580 55804 97636 55860
rect 97804 55916 97860 55972
rect 95564 54236 95620 54292
rect 95340 52108 95396 52164
rect 95452 50092 95508 50148
rect 96636 54122 96692 54124
rect 96636 54070 96638 54122
rect 96638 54070 96690 54122
rect 96690 54070 96692 54122
rect 96636 54068 96692 54070
rect 96740 54122 96796 54124
rect 96740 54070 96742 54122
rect 96742 54070 96794 54122
rect 96794 54070 96796 54122
rect 96740 54068 96796 54070
rect 96844 54122 96900 54124
rect 96844 54070 96846 54122
rect 96846 54070 96898 54122
rect 96898 54070 96900 54122
rect 96844 54068 96900 54070
rect 97692 53730 97748 53732
rect 97692 53678 97694 53730
rect 97694 53678 97746 53730
rect 97746 53678 97748 53730
rect 97692 53676 97748 53678
rect 95676 53170 95732 53172
rect 95676 53118 95678 53170
rect 95678 53118 95730 53170
rect 95730 53118 95732 53170
rect 95676 53116 95732 53118
rect 96908 53116 96964 53172
rect 96124 52946 96180 52948
rect 96124 52894 96126 52946
rect 96126 52894 96178 52946
rect 96178 52894 96180 52946
rect 96124 52892 96180 52894
rect 96124 52556 96180 52612
rect 95452 49922 95508 49924
rect 95452 49870 95454 49922
rect 95454 49870 95506 49922
rect 95506 49870 95508 49922
rect 95452 49868 95508 49870
rect 95228 48860 95284 48916
rect 95340 49644 95396 49700
rect 94892 47740 94948 47796
rect 94556 47180 94612 47236
rect 95228 47346 95284 47348
rect 95228 47294 95230 47346
rect 95230 47294 95282 47346
rect 95282 47294 95284 47346
rect 95228 47292 95284 47294
rect 95116 46396 95172 46452
rect 96236 51884 96292 51940
rect 96236 51490 96292 51492
rect 96236 51438 96238 51490
rect 96238 51438 96290 51490
rect 96290 51438 96292 51490
rect 96236 51436 96292 51438
rect 96348 50316 96404 50372
rect 95676 49980 95732 50036
rect 96124 50034 96180 50036
rect 96124 49982 96126 50034
rect 96126 49982 96178 50034
rect 96178 49982 96180 50034
rect 96124 49980 96180 49982
rect 95788 49922 95844 49924
rect 95788 49870 95790 49922
rect 95790 49870 95842 49922
rect 95842 49870 95844 49922
rect 95788 49868 95844 49870
rect 95564 47404 95620 47460
rect 95564 46844 95620 46900
rect 95676 49756 95732 49812
rect 96636 52554 96692 52556
rect 96636 52502 96638 52554
rect 96638 52502 96690 52554
rect 96690 52502 96692 52554
rect 96636 52500 96692 52502
rect 96740 52554 96796 52556
rect 96740 52502 96742 52554
rect 96742 52502 96794 52554
rect 96794 52502 96796 52554
rect 96740 52500 96796 52502
rect 96844 52554 96900 52556
rect 96844 52502 96846 52554
rect 96846 52502 96898 52554
rect 96898 52502 96900 52554
rect 96844 52500 96900 52502
rect 97580 52946 97636 52948
rect 97580 52894 97582 52946
rect 97582 52894 97634 52946
rect 97634 52894 97636 52946
rect 97580 52892 97636 52894
rect 97132 52834 97188 52836
rect 97132 52782 97134 52834
rect 97134 52782 97186 52834
rect 97186 52782 97188 52834
rect 97132 52780 97188 52782
rect 98028 53676 98084 53732
rect 97468 51548 97524 51604
rect 97692 51436 97748 51492
rect 96636 50986 96692 50988
rect 96636 50934 96638 50986
rect 96638 50934 96690 50986
rect 96690 50934 96692 50986
rect 96636 50932 96692 50934
rect 96740 50986 96796 50988
rect 96740 50934 96742 50986
rect 96742 50934 96794 50986
rect 96794 50934 96796 50986
rect 96740 50932 96796 50934
rect 96844 50986 96900 50988
rect 96844 50934 96846 50986
rect 96846 50934 96898 50986
rect 96898 50934 96900 50986
rect 96844 50932 96900 50934
rect 97468 50092 97524 50148
rect 97356 49922 97412 49924
rect 97356 49870 97358 49922
rect 97358 49870 97410 49922
rect 97410 49870 97412 49922
rect 97356 49868 97412 49870
rect 96636 49418 96692 49420
rect 96636 49366 96638 49418
rect 96638 49366 96690 49418
rect 96690 49366 96692 49418
rect 96636 49364 96692 49366
rect 96740 49418 96796 49420
rect 96740 49366 96742 49418
rect 96742 49366 96794 49418
rect 96794 49366 96796 49418
rect 96740 49364 96796 49366
rect 96844 49418 96900 49420
rect 96844 49366 96846 49418
rect 96846 49366 96898 49418
rect 96898 49366 96900 49418
rect 96844 49364 96900 49366
rect 96236 48300 96292 48356
rect 97468 48354 97524 48356
rect 97468 48302 97470 48354
rect 97470 48302 97522 48354
rect 97522 48302 97524 48354
rect 97468 48300 97524 48302
rect 97244 48076 97300 48132
rect 96636 47850 96692 47852
rect 96236 47740 96292 47796
rect 96636 47798 96638 47850
rect 96638 47798 96690 47850
rect 96690 47798 96692 47850
rect 96636 47796 96692 47798
rect 96740 47850 96796 47852
rect 96740 47798 96742 47850
rect 96742 47798 96794 47850
rect 96794 47798 96796 47850
rect 96740 47796 96796 47798
rect 96844 47850 96900 47852
rect 96844 47798 96846 47850
rect 96846 47798 96898 47850
rect 96898 47798 96900 47850
rect 96844 47796 96900 47798
rect 96460 47458 96516 47460
rect 96460 47406 96462 47458
rect 96462 47406 96514 47458
rect 96514 47406 96516 47458
rect 96460 47404 96516 47406
rect 96012 46898 96068 46900
rect 96012 46846 96014 46898
rect 96014 46846 96066 46898
rect 96066 46846 96068 46898
rect 96012 46844 96068 46846
rect 96796 47068 96852 47124
rect 97804 51884 97860 51940
rect 97916 49810 97972 49812
rect 97916 49758 97918 49810
rect 97918 49758 97970 49810
rect 97970 49758 97972 49810
rect 97916 49756 97972 49758
rect 97580 47404 97636 47460
rect 97356 46396 97412 46452
rect 96636 46282 96692 46284
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 94332 42866 94388 42868
rect 94332 42814 94334 42866
rect 94334 42814 94386 42866
rect 94386 42814 94388 42866
rect 94332 42812 94388 42814
rect 94556 42812 94612 42868
rect 94332 41858 94388 41860
rect 94332 41806 94334 41858
rect 94334 41806 94386 41858
rect 94386 41806 94388 41858
rect 94332 41804 94388 41806
rect 93996 40460 94052 40516
rect 93100 38780 93156 38836
rect 94220 38780 94276 38836
rect 93884 38556 93940 38612
rect 93100 37378 93156 37380
rect 93100 37326 93102 37378
rect 93102 37326 93154 37378
rect 93154 37326 93156 37378
rect 93100 37324 93156 37326
rect 94108 37938 94164 37940
rect 94108 37886 94110 37938
rect 94110 37886 94162 37938
rect 94162 37886 94164 37938
rect 94108 37884 94164 37886
rect 94332 38556 94388 38612
rect 95788 44380 95844 44436
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 95900 43820 95956 43876
rect 95564 43650 95620 43652
rect 95564 43598 95566 43650
rect 95566 43598 95618 43650
rect 95618 43598 95620 43650
rect 95564 43596 95620 43598
rect 95564 42812 95620 42868
rect 95788 43708 95844 43764
rect 95004 42476 95060 42532
rect 95340 42476 95396 42532
rect 94892 41692 94948 41748
rect 95228 41970 95284 41972
rect 95228 41918 95230 41970
rect 95230 41918 95282 41970
rect 95282 41918 95284 41970
rect 95228 41916 95284 41918
rect 94892 39730 94948 39732
rect 94892 39678 94894 39730
rect 94894 39678 94946 39730
rect 94946 39678 94948 39730
rect 94892 39676 94948 39678
rect 96236 43708 96292 43764
rect 97020 43708 97076 43764
rect 98252 47964 98308 48020
rect 97692 43596 97748 43652
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 95676 41804 95732 41860
rect 96124 42812 96180 42868
rect 95340 41298 95396 41300
rect 95340 41246 95342 41298
rect 95342 41246 95394 41298
rect 95394 41246 95396 41298
rect 95340 41244 95396 41246
rect 96012 41746 96068 41748
rect 96012 41694 96014 41746
rect 96014 41694 96066 41746
rect 96066 41694 96068 41746
rect 96012 41692 96068 41694
rect 95340 39676 95396 39732
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 96796 41074 96852 41076
rect 96796 41022 96798 41074
rect 96798 41022 96850 41074
rect 96850 41022 96852 41074
rect 96796 41020 96852 41022
rect 96348 40572 96404 40628
rect 96124 40514 96180 40516
rect 96124 40462 96126 40514
rect 96126 40462 96178 40514
rect 96178 40462 96180 40514
rect 96124 40460 96180 40462
rect 97356 41132 97412 41188
rect 96908 40460 96964 40516
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 97580 41186 97636 41188
rect 97580 41134 97582 41186
rect 97582 41134 97634 41186
rect 97634 41134 97636 41186
rect 97580 41132 97636 41134
rect 97468 40572 97524 40628
rect 96460 38780 96516 38836
rect 95788 38668 95844 38724
rect 95452 38556 95508 38612
rect 96236 38556 96292 38612
rect 95452 37938 95508 37940
rect 95452 37886 95454 37938
rect 95454 37886 95506 37938
rect 95506 37886 95508 37938
rect 95452 37884 95508 37886
rect 93772 36652 93828 36708
rect 95228 36706 95284 36708
rect 95228 36654 95230 36706
rect 95230 36654 95282 36706
rect 95282 36654 95284 36706
rect 95228 36652 95284 36654
rect 93212 36594 93268 36596
rect 93212 36542 93214 36594
rect 93214 36542 93266 36594
rect 93266 36542 93268 36594
rect 93212 36540 93268 36542
rect 93772 36482 93828 36484
rect 93772 36430 93774 36482
rect 93774 36430 93826 36482
rect 93826 36430 93828 36482
rect 93772 36428 93828 36430
rect 92876 35196 92932 35252
rect 93660 34412 93716 34468
rect 93996 34412 94052 34468
rect 92428 34076 92484 34132
rect 90748 33964 90804 34020
rect 90188 33628 90244 33684
rect 92204 34018 92260 34020
rect 92204 33966 92206 34018
rect 92206 33966 92258 34018
rect 92258 33966 92260 34018
rect 92204 33964 92260 33966
rect 91644 33628 91700 33684
rect 93100 34242 93156 34244
rect 93100 34190 93102 34242
rect 93102 34190 93154 34242
rect 93154 34190 93156 34242
rect 93100 34188 93156 34190
rect 92764 33628 92820 33684
rect 92428 33346 92484 33348
rect 92428 33294 92430 33346
rect 92430 33294 92482 33346
rect 92482 33294 92484 33346
rect 92428 33292 92484 33294
rect 95564 37212 95620 37268
rect 96012 37266 96068 37268
rect 96012 37214 96014 37266
rect 96014 37214 96066 37266
rect 96066 37214 96068 37266
rect 96012 37212 96068 37214
rect 95452 36540 95508 36596
rect 95788 36540 95844 36596
rect 95340 36428 95396 36484
rect 98028 41970 98084 41972
rect 98028 41918 98030 41970
rect 98030 41918 98082 41970
rect 98082 41918 98084 41970
rect 98028 41916 98084 41918
rect 97468 38780 97524 38836
rect 97020 38668 97076 38724
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 94332 34300 94388 34356
rect 96124 35196 96180 35252
rect 93996 33516 94052 33572
rect 95228 34354 95284 34356
rect 95228 34302 95230 34354
rect 95230 34302 95282 34354
rect 95282 34302 95284 34354
rect 95228 34300 95284 34302
rect 96124 34300 96180 34356
rect 95564 34130 95620 34132
rect 95564 34078 95566 34130
rect 95566 34078 95618 34130
rect 95618 34078 95620 34130
rect 95564 34076 95620 34078
rect 94444 33292 94500 33348
rect 94668 32786 94724 32788
rect 94668 32734 94670 32786
rect 94670 32734 94722 32786
rect 94722 32734 94724 32786
rect 94668 32732 94724 32734
rect 90972 32562 91028 32564
rect 90972 32510 90974 32562
rect 90974 32510 91026 32562
rect 91026 32510 91028 32562
rect 90972 32508 91028 32510
rect 91532 32562 91588 32564
rect 91532 32510 91534 32562
rect 91534 32510 91586 32562
rect 91586 32510 91588 32562
rect 91532 32508 91588 32510
rect 95788 33516 95844 33572
rect 98028 38722 98084 38724
rect 98028 38670 98030 38722
rect 98030 38670 98082 38722
rect 98082 38670 98084 38722
rect 98028 38668 98084 38670
rect 98252 39676 98308 39732
rect 98140 38556 98196 38612
rect 97580 37212 97636 37268
rect 97132 36540 97188 36596
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 97132 34354 97188 34356
rect 97132 34302 97134 34354
rect 97134 34302 97186 34354
rect 97186 34302 97188 34354
rect 97132 34300 97188 34302
rect 97244 34076 97300 34132
rect 97468 34300 97524 34356
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 96236 32732 96292 32788
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 90748 31836 90804 31892
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 94892 25282 94948 25284
rect 94892 25230 94894 25282
rect 94894 25230 94946 25282
rect 94946 25230 94948 25282
rect 94892 25228 94948 25230
rect 95228 25228 95284 25284
rect 95788 25282 95844 25284
rect 95788 25230 95790 25282
rect 95790 25230 95842 25282
rect 95842 25230 95844 25282
rect 95788 25228 95844 25230
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 93436 3388 93492 3444
rect 89628 3276 89684 3332
rect 82460 2940 82516 2996
rect 93996 3442 94052 3444
rect 93996 3390 93998 3442
rect 93998 3390 94050 3442
rect 94050 3390 94052 3442
rect 93996 3388 94052 3390
rect 93660 2828 93716 2884
<< metal3 >>
rect 4466 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4750 96460
rect 35186 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35470 96460
rect 65906 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66190 96460
rect 96626 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96910 96460
rect 93426 96124 93436 96180
rect 93492 96124 94332 96180
rect 94388 96124 94398 96180
rect 7858 96012 7868 96068
rect 7924 96012 8316 96068
rect 8372 96012 47964 96068
rect 48020 96012 48030 96068
rect 93090 96012 93100 96068
rect 93156 96012 93884 96068
rect 93940 96012 97468 96068
rect 97524 96012 97534 96068
rect 20290 95788 20300 95844
rect 20356 95788 21308 95844
rect 21364 95788 27692 95844
rect 27748 95788 27758 95844
rect 70018 95788 70028 95844
rect 70084 95788 70476 95844
rect 70532 95788 77980 95844
rect 78036 95788 78046 95844
rect 19826 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20110 95676
rect 50546 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50830 95676
rect 81266 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81550 95676
rect 4466 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4750 94892
rect 35186 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35470 94892
rect 65906 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66190 94892
rect 96626 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96910 94892
rect 19826 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20110 94108
rect 50546 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50830 94108
rect 81266 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81550 94108
rect 4466 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4750 93324
rect 35186 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35470 93324
rect 65906 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66190 93324
rect 96626 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96910 93324
rect 19826 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20110 92540
rect 50546 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50830 92540
rect 81266 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81550 92540
rect 4466 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4750 91756
rect 35186 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35470 91756
rect 65906 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66190 91756
rect 96626 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96910 91756
rect 19826 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20110 90972
rect 50546 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50830 90972
rect 81266 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81550 90972
rect 4466 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4750 90188
rect 35186 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35470 90188
rect 65906 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66190 90188
rect 96626 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96910 90188
rect 19826 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20110 89404
rect 50546 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50830 89404
rect 81266 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81550 89404
rect 70466 88844 70476 88900
rect 70532 88844 71596 88900
rect 71652 88844 71662 88900
rect 4466 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4750 88620
rect 35186 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35470 88620
rect 65906 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66190 88620
rect 96626 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96910 88620
rect 3266 88284 3276 88340
rect 3332 88284 12572 88340
rect 12628 88284 12638 88340
rect 59042 87836 59052 87892
rect 59108 87836 59612 87892
rect 59668 87836 60284 87892
rect 60340 87836 62524 87892
rect 62580 87836 64428 87892
rect 64484 87836 71932 87892
rect 71988 87836 71998 87892
rect 19826 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20110 87836
rect 50546 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50830 87836
rect 81266 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81550 87836
rect 62738 87500 62748 87556
rect 62804 87500 64316 87556
rect 64372 87500 64382 87556
rect 88386 87500 88396 87556
rect 88452 87500 89516 87556
rect 89572 87500 90860 87556
rect 90916 87500 90926 87556
rect 0 87444 800 87472
rect 0 87388 1708 87444
rect 1764 87388 1774 87444
rect 71922 87388 71932 87444
rect 71988 87388 73164 87444
rect 73220 87388 73230 87444
rect 92642 87388 92652 87444
rect 92708 87388 94556 87444
rect 94612 87388 95116 87444
rect 95172 87388 95182 87444
rect 0 87360 800 87388
rect 54226 87276 54236 87332
rect 54292 87276 54796 87332
rect 54852 87276 55020 87332
rect 55076 87276 55086 87332
rect 60498 87276 60508 87332
rect 60564 87276 61852 87332
rect 61908 87276 61918 87332
rect 67442 87276 67452 87332
rect 67508 87276 68236 87332
rect 68292 87276 68302 87332
rect 72482 87276 72492 87332
rect 72548 87276 73724 87332
rect 73780 87276 73790 87332
rect 53554 87164 53564 87220
rect 53620 87164 56028 87220
rect 56084 87164 57484 87220
rect 57540 87164 57820 87220
rect 57876 87164 58380 87220
rect 58436 87164 58446 87220
rect 62402 87164 62412 87220
rect 62468 87164 63084 87220
rect 63140 87164 63756 87220
rect 63812 87164 63822 87220
rect 4466 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4750 87052
rect 35186 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35470 87052
rect 65906 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66190 87052
rect 96626 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96910 87052
rect 57586 86940 57596 86996
rect 57652 86940 60844 86996
rect 60900 86940 60910 86996
rect 87042 86828 87052 86884
rect 87108 86828 87612 86884
rect 87668 86828 87678 86884
rect 56466 86716 56476 86772
rect 56532 86716 57596 86772
rect 57652 86716 59948 86772
rect 60004 86716 60620 86772
rect 60676 86716 62188 86772
rect 62244 86716 63308 86772
rect 63364 86716 63374 86772
rect 69234 86604 69244 86660
rect 69300 86604 69804 86660
rect 69860 86604 69870 86660
rect 70242 86604 70252 86660
rect 70308 86604 71708 86660
rect 71764 86604 71774 86660
rect 73378 86604 73388 86660
rect 73444 86604 73724 86660
rect 73780 86604 74396 86660
rect 74452 86604 75516 86660
rect 75572 86604 75582 86660
rect 68562 86492 68572 86548
rect 68628 86492 71372 86548
rect 71428 86492 71438 86548
rect 74946 86492 74956 86548
rect 75012 86492 75740 86548
rect 75796 86492 75806 86548
rect 85586 86492 85596 86548
rect 85652 86492 88732 86548
rect 88788 86492 89740 86548
rect 89796 86492 89806 86548
rect 65538 86380 65548 86436
rect 65604 86380 66668 86436
rect 66724 86380 66734 86436
rect 68338 86380 68348 86436
rect 68404 86380 69468 86436
rect 69524 86380 69534 86436
rect 70354 86380 70364 86436
rect 70420 86380 70588 86436
rect 70644 86380 71036 86436
rect 71092 86380 71102 86436
rect 81218 86380 81228 86436
rect 81284 86380 81900 86436
rect 81956 86380 82460 86436
rect 82516 86380 83132 86436
rect 83188 86380 83198 86436
rect 87042 86380 87052 86436
rect 87108 86380 88172 86436
rect 88228 86380 89180 86436
rect 89236 86380 89246 86436
rect 58706 86268 58716 86324
rect 58772 86268 59276 86324
rect 59332 86268 59342 86324
rect 64530 86268 64540 86324
rect 64596 86268 65772 86324
rect 65828 86268 65838 86324
rect 67172 86268 70140 86324
rect 70196 86268 70700 86324
rect 70756 86268 71932 86324
rect 71988 86268 71998 86324
rect 87938 86268 87948 86324
rect 88004 86268 89292 86324
rect 89348 86268 91532 86324
rect 91588 86268 91598 86324
rect 19826 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20110 86268
rect 50546 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50830 86268
rect 61506 86156 61516 86212
rect 61572 86156 63420 86212
rect 63476 86156 63486 86212
rect 67172 86100 67228 86268
rect 81266 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81550 86268
rect 54674 86044 54684 86100
rect 54740 86044 56476 86100
rect 56532 86044 57708 86100
rect 57764 86044 67228 86100
rect 70354 86044 70364 86100
rect 70420 86044 71596 86100
rect 71652 86044 71662 86100
rect 72706 86044 72716 86100
rect 72772 86044 73388 86100
rect 73444 86044 73454 86100
rect 77858 86044 77868 86100
rect 77924 86044 79212 86100
rect 79268 86044 79278 86100
rect 54002 85932 54012 85988
rect 54068 85932 55692 85988
rect 55748 85932 56700 85988
rect 56756 85932 56766 85988
rect 58258 85932 58268 85988
rect 58324 85932 59836 85988
rect 59892 85932 59902 85988
rect 87266 85932 87276 85988
rect 87332 85932 87724 85988
rect 87780 85932 87790 85988
rect 61730 85820 61740 85876
rect 61796 85820 63084 85876
rect 63140 85820 63150 85876
rect 65762 85820 65772 85876
rect 65828 85820 67228 85876
rect 67284 85820 67294 85876
rect 75292 85820 76524 85876
rect 76580 85820 76590 85876
rect 75292 85764 75348 85820
rect 55794 85708 55804 85764
rect 55860 85708 60508 85764
rect 60564 85708 60574 85764
rect 60946 85708 60956 85764
rect 61012 85708 62412 85764
rect 62468 85708 62478 85764
rect 62962 85708 62972 85764
rect 63028 85708 63868 85764
rect 63924 85708 64316 85764
rect 64372 85708 65436 85764
rect 65492 85708 65502 85764
rect 67442 85708 67452 85764
rect 67508 85708 69468 85764
rect 69524 85708 70476 85764
rect 70532 85708 70542 85764
rect 74722 85708 74732 85764
rect 74788 85708 75292 85764
rect 75348 85708 75358 85764
rect 76066 85708 76076 85764
rect 76132 85708 77420 85764
rect 77476 85708 78204 85764
rect 78260 85708 78270 85764
rect 78866 85708 78876 85764
rect 78932 85708 79660 85764
rect 79716 85708 79726 85764
rect 82338 85708 82348 85764
rect 82404 85708 88060 85764
rect 88116 85708 88126 85764
rect 70476 85652 70532 85708
rect 70476 85596 73164 85652
rect 73220 85596 73230 85652
rect 79762 85596 79772 85652
rect 79828 85596 80444 85652
rect 80500 85596 80510 85652
rect 81666 85596 81676 85652
rect 81732 85596 82796 85652
rect 82852 85596 82862 85652
rect 4466 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4750 85484
rect 35186 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35470 85484
rect 65906 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66190 85484
rect 96626 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96910 85484
rect 59378 85260 59388 85316
rect 59444 85260 60396 85316
rect 60452 85260 60462 85316
rect 86482 85260 86492 85316
rect 86548 85260 88844 85316
rect 88900 85260 88910 85316
rect 56578 85148 56588 85204
rect 56644 85148 57260 85204
rect 57316 85148 59500 85204
rect 59556 85148 59566 85204
rect 87490 85148 87500 85204
rect 87556 85148 88172 85204
rect 88228 85148 89180 85204
rect 89236 85148 89246 85204
rect 93538 85148 93548 85204
rect 93604 85148 94892 85204
rect 94948 85148 94958 85204
rect 82562 85036 82572 85092
rect 82628 85036 83468 85092
rect 83524 85036 83534 85092
rect 91186 85036 91196 85092
rect 91252 85036 93436 85092
rect 93492 85036 93502 85092
rect 67106 84924 67116 84980
rect 67172 84924 67340 84980
rect 67396 84924 74844 84980
rect 74900 84924 75628 84980
rect 75684 84924 75694 84980
rect 92306 84924 92316 84980
rect 92372 84924 93772 84980
rect 93828 84924 93838 84980
rect 53778 84812 53788 84868
rect 53844 84812 54460 84868
rect 54516 84812 54526 84868
rect 63746 84812 63756 84868
rect 63812 84812 66220 84868
rect 66276 84812 66286 84868
rect 19826 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20110 84700
rect 50546 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50830 84700
rect 81266 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81550 84700
rect 65762 84476 65772 84532
rect 65828 84476 66556 84532
rect 66612 84476 66622 84532
rect 73938 84476 73948 84532
rect 74004 84476 90524 84532
rect 90580 84476 92204 84532
rect 92260 84476 92270 84532
rect 94434 84476 94444 84532
rect 94500 84476 95564 84532
rect 95620 84476 95630 84532
rect 67106 84364 67116 84420
rect 67172 84364 68012 84420
rect 68068 84364 68078 84420
rect 81666 84364 81676 84420
rect 81732 84364 84924 84420
rect 84980 84364 84990 84420
rect 87714 84364 87724 84420
rect 87780 84364 89292 84420
rect 89348 84364 89358 84420
rect 96338 84364 96348 84420
rect 96404 84364 97804 84420
rect 97860 84364 97870 84420
rect 56914 84252 56924 84308
rect 56980 84252 58828 84308
rect 58884 84252 64316 84308
rect 64372 84252 66444 84308
rect 66500 84252 66510 84308
rect 73602 84252 73612 84308
rect 73668 84252 74620 84308
rect 74676 84252 75516 84308
rect 75572 84252 77420 84308
rect 77476 84252 78764 84308
rect 78820 84252 79548 84308
rect 79604 84252 80444 84308
rect 80500 84252 81452 84308
rect 81508 84252 83020 84308
rect 83076 84252 83086 84308
rect 88498 84252 88508 84308
rect 88564 84252 90188 84308
rect 90244 84252 90254 84308
rect 55794 84140 55804 84196
rect 55860 84140 56476 84196
rect 56532 84140 57372 84196
rect 57428 84140 57438 84196
rect 80546 84140 80556 84196
rect 80612 84140 82124 84196
rect 82180 84140 82190 84196
rect 89394 84140 89404 84196
rect 89460 84140 91532 84196
rect 91588 84140 94220 84196
rect 94276 84140 94286 84196
rect 64418 84028 64428 84084
rect 64484 84028 65100 84084
rect 65156 84028 67340 84084
rect 67396 84028 67676 84084
rect 67732 84028 67742 84084
rect 75394 84028 75404 84084
rect 75460 84028 76412 84084
rect 76468 84028 77420 84084
rect 77476 84028 77486 84084
rect 82674 84028 82684 84084
rect 82740 84028 84924 84084
rect 84980 84028 84990 84084
rect 88274 84028 88284 84084
rect 88340 84028 89516 84084
rect 89572 84028 89582 84084
rect 4466 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4750 83916
rect 35186 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35470 83916
rect 65906 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66190 83916
rect 96626 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96910 83916
rect 85586 83692 85596 83748
rect 85652 83692 87388 83748
rect 87444 83692 88620 83748
rect 88676 83692 88686 83748
rect 53218 83580 53228 83636
rect 53284 83580 53676 83636
rect 53732 83580 54460 83636
rect 54516 83580 54526 83636
rect 94322 83580 94332 83636
rect 94388 83580 95788 83636
rect 95844 83580 95854 83636
rect 88386 83468 88396 83524
rect 88452 83468 90748 83524
rect 90804 83468 91532 83524
rect 91588 83468 91598 83524
rect 92194 83468 92204 83524
rect 92260 83468 96236 83524
rect 96292 83468 96302 83524
rect 76402 83356 76412 83412
rect 76468 83356 78540 83412
rect 78596 83356 78606 83412
rect 80434 83356 80444 83412
rect 80500 83356 82012 83412
rect 82068 83356 83580 83412
rect 83636 83356 83646 83412
rect 52434 83244 52444 83300
rect 52500 83244 54124 83300
rect 54180 83244 54190 83300
rect 71250 83244 71260 83300
rect 71316 83244 71596 83300
rect 71652 83244 73164 83300
rect 73220 83244 87612 83300
rect 87668 83244 88844 83300
rect 88900 83244 89628 83300
rect 89684 83244 89694 83300
rect 19826 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20110 83132
rect 50546 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50830 83132
rect 81266 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81550 83132
rect 52210 82684 52220 82740
rect 52276 82684 52892 82740
rect 52948 82684 56924 82740
rect 56980 82684 56990 82740
rect 83906 82684 83916 82740
rect 83972 82684 85036 82740
rect 85092 82684 85102 82740
rect 58930 82572 58940 82628
rect 58996 82572 60396 82628
rect 60452 82572 60462 82628
rect 73266 82572 73276 82628
rect 73332 82572 73836 82628
rect 73892 82572 74956 82628
rect 75012 82572 75022 82628
rect 82002 82572 82012 82628
rect 82068 82572 85260 82628
rect 85316 82572 86604 82628
rect 86660 82572 87612 82628
rect 87668 82572 90412 82628
rect 90468 82572 90478 82628
rect 4466 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4750 82348
rect 35186 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35470 82348
rect 65906 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66190 82348
rect 96626 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96910 82348
rect 54114 82236 54124 82292
rect 54180 82236 54908 82292
rect 54964 82236 54974 82292
rect 68674 82236 68684 82292
rect 68740 82236 69244 82292
rect 69300 82236 69310 82292
rect 77522 82236 77532 82292
rect 77588 82236 79212 82292
rect 79268 82236 80444 82292
rect 80500 82236 80510 82292
rect 80658 82236 80668 82292
rect 80724 82236 81452 82292
rect 81508 82236 83020 82292
rect 83076 82236 83086 82292
rect 83458 82236 83468 82292
rect 83524 82236 84140 82292
rect 84196 82236 84206 82292
rect 78932 82124 95788 82180
rect 95844 82124 95854 82180
rect 78932 82068 78988 82124
rect 52658 82012 52668 82068
rect 52724 82012 53564 82068
rect 53620 82012 53630 82068
rect 60834 82012 60844 82068
rect 60900 82012 63980 82068
rect 64036 82012 64046 82068
rect 75394 82012 75404 82068
rect 75460 82012 77532 82068
rect 77588 82012 77598 82068
rect 77858 82012 77868 82068
rect 77924 82012 78652 82068
rect 78708 82012 78988 82068
rect 94098 82012 94108 82068
rect 94164 82012 97356 82068
rect 97412 82012 97422 82068
rect 52770 81900 52780 81956
rect 52836 81900 53340 81956
rect 53396 81900 54124 81956
rect 54180 81900 54190 81956
rect 62178 81900 62188 81956
rect 62244 81900 62524 81956
rect 62580 81900 63644 81956
rect 63700 81900 63710 81956
rect 80322 81900 80332 81956
rect 80388 81900 82684 81956
rect 82740 81900 82750 81956
rect 72818 81788 72828 81844
rect 72884 81788 73612 81844
rect 73668 81788 73892 81844
rect 73836 81732 73892 81788
rect 55010 81676 55020 81732
rect 55076 81676 56588 81732
rect 56644 81676 56654 81732
rect 59714 81676 59724 81732
rect 59780 81676 60284 81732
rect 60340 81676 63420 81732
rect 63476 81676 64092 81732
rect 64148 81676 64428 81732
rect 64484 81676 73276 81732
rect 73332 81676 73342 81732
rect 73826 81676 73836 81732
rect 73892 81676 74284 81732
rect 74340 81676 74844 81732
rect 74900 81676 74910 81732
rect 75730 81676 75740 81732
rect 75796 81676 76524 81732
rect 76580 81676 77196 81732
rect 77252 81676 77262 81732
rect 83682 81676 83692 81732
rect 83748 81676 84812 81732
rect 84868 81676 84878 81732
rect 92418 81676 92428 81732
rect 92484 81676 93884 81732
rect 93940 81676 93950 81732
rect 82898 81564 82908 81620
rect 82964 81564 84252 81620
rect 84308 81564 85260 81620
rect 85316 81564 85326 81620
rect 19826 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20110 81564
rect 50546 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50830 81564
rect 81266 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81550 81564
rect 78932 81452 80556 81508
rect 80612 81452 80622 81508
rect 78932 81396 78988 81452
rect 65762 81340 65772 81396
rect 65828 81340 66332 81396
rect 66388 81340 69468 81396
rect 69524 81340 69692 81396
rect 69748 81340 69758 81396
rect 73826 81340 73836 81396
rect 73892 81340 75068 81396
rect 75124 81340 75292 81396
rect 75348 81340 78988 81396
rect 80434 81340 80444 81396
rect 80500 81340 90748 81396
rect 90692 81284 90748 81340
rect 50306 81228 50316 81284
rect 50372 81228 54012 81284
rect 54068 81228 54078 81284
rect 80108 81228 80668 81284
rect 80724 81228 80734 81284
rect 81666 81228 81676 81284
rect 81732 81228 82348 81284
rect 82404 81228 82414 81284
rect 90692 81228 92204 81284
rect 92260 81228 92270 81284
rect 80108 81172 80164 81228
rect 49746 81116 49756 81172
rect 49812 81116 51212 81172
rect 51268 81116 51660 81172
rect 51716 81116 53340 81172
rect 53396 81116 53406 81172
rect 71474 81116 71484 81172
rect 71540 81116 80108 81172
rect 80164 81116 80174 81172
rect 80434 81116 80444 81172
rect 80500 81116 81564 81172
rect 81620 81116 82124 81172
rect 82180 81116 82190 81172
rect 68114 81004 68124 81060
rect 68180 81004 70140 81060
rect 70196 81004 70206 81060
rect 80546 81004 80556 81060
rect 80612 81004 82460 81060
rect 82516 81004 82526 81060
rect 83682 81004 83692 81060
rect 83748 81004 84364 81060
rect 84420 81004 84588 81060
rect 84644 81004 84654 81060
rect 93202 81004 93212 81060
rect 93268 81004 94668 81060
rect 94724 81004 94734 81060
rect 95554 81004 95564 81060
rect 95620 81004 97244 81060
rect 97300 81004 97310 81060
rect 51090 80892 51100 80948
rect 51156 80892 53452 80948
rect 53508 80892 55020 80948
rect 55076 80892 55086 80948
rect 69682 80892 69692 80948
rect 69748 80892 70588 80948
rect 70644 80892 71708 80948
rect 71764 80892 71774 80948
rect 79538 80892 79548 80948
rect 79604 80892 81452 80948
rect 81508 80892 81518 80948
rect 80322 80780 80332 80836
rect 80388 80780 82908 80836
rect 82964 80780 82974 80836
rect 4466 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4750 80780
rect 35186 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35470 80780
rect 65906 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66190 80780
rect 96626 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96910 80780
rect 63634 80668 63644 80724
rect 63700 80668 64204 80724
rect 64260 80668 64270 80724
rect 74722 80668 74732 80724
rect 74788 80668 74798 80724
rect 78306 80668 78316 80724
rect 78372 80668 79324 80724
rect 79380 80668 79390 80724
rect 82002 80668 82012 80724
rect 82068 80668 84140 80724
rect 84196 80668 86716 80724
rect 86772 80668 90972 80724
rect 91028 80668 91196 80724
rect 91252 80668 92428 80724
rect 92484 80668 93100 80724
rect 93156 80668 93166 80724
rect 93538 80668 93548 80724
rect 93604 80668 93884 80724
rect 93940 80668 94556 80724
rect 94612 80668 94622 80724
rect 74732 80612 74788 80668
rect 56018 80556 56028 80612
rect 56084 80556 56924 80612
rect 56980 80556 56990 80612
rect 61506 80556 61516 80612
rect 61572 80556 62636 80612
rect 62692 80556 63420 80612
rect 63476 80556 63486 80612
rect 69234 80556 69244 80612
rect 69300 80556 70476 80612
rect 70532 80556 70542 80612
rect 74732 80556 75964 80612
rect 76020 80556 76030 80612
rect 81106 80556 81116 80612
rect 81172 80556 83580 80612
rect 83636 80556 83646 80612
rect 95442 80556 95452 80612
rect 95508 80556 96124 80612
rect 96180 80556 97804 80612
rect 97860 80556 97870 80612
rect 54226 80444 54236 80500
rect 54292 80444 54908 80500
rect 54964 80444 54974 80500
rect 56354 80444 56364 80500
rect 56420 80444 57036 80500
rect 57092 80444 57484 80500
rect 57540 80444 57550 80500
rect 61394 80444 61404 80500
rect 61460 80444 62972 80500
rect 63028 80444 63038 80500
rect 67172 80444 70700 80500
rect 70756 80444 70766 80500
rect 74498 80444 74508 80500
rect 74564 80444 75180 80500
rect 75236 80444 75246 80500
rect 86034 80444 86044 80500
rect 86100 80444 86828 80500
rect 86884 80444 86894 80500
rect 95330 80444 95340 80500
rect 95396 80444 97692 80500
rect 97748 80444 97758 80500
rect 67172 80388 67228 80444
rect 55346 80332 55356 80388
rect 55412 80332 56812 80388
rect 56868 80332 56878 80388
rect 57138 80332 57148 80388
rect 57204 80332 57372 80388
rect 57428 80332 57596 80388
rect 57652 80332 67228 80388
rect 68002 80332 68012 80388
rect 68068 80332 70028 80388
rect 70084 80332 70094 80388
rect 70354 80332 70364 80388
rect 70420 80332 71372 80388
rect 71428 80332 71438 80388
rect 82898 80332 82908 80388
rect 82964 80332 84252 80388
rect 84308 80332 85372 80388
rect 85428 80332 85596 80388
rect 85652 80332 85662 80388
rect 93314 80332 93324 80388
rect 93380 80332 94892 80388
rect 94948 80332 94958 80388
rect 57148 80276 57204 80332
rect 56130 80220 56140 80276
rect 56196 80220 57204 80276
rect 68562 80220 68572 80276
rect 68628 80220 69468 80276
rect 69524 80220 69534 80276
rect 70802 80220 70812 80276
rect 70868 80220 71484 80276
rect 71540 80220 78988 80276
rect 81330 80220 81340 80276
rect 81396 80220 83020 80276
rect 83076 80220 83086 80276
rect 83570 80220 83580 80276
rect 83636 80220 84476 80276
rect 84532 80220 84700 80276
rect 84756 80220 84766 80276
rect 94322 80220 94332 80276
rect 94388 80220 95788 80276
rect 95844 80220 95854 80276
rect 78932 80164 78988 80220
rect 53218 80108 53228 80164
rect 53284 80108 55468 80164
rect 68226 80108 68236 80164
rect 68292 80108 69244 80164
rect 69300 80108 70140 80164
rect 70196 80108 70206 80164
rect 70354 80108 70364 80164
rect 70420 80108 71708 80164
rect 71764 80108 73836 80164
rect 73892 80108 76188 80164
rect 76244 80108 76254 80164
rect 78932 80108 82068 80164
rect 82226 80108 82236 80164
rect 82292 80108 83244 80164
rect 83300 80108 83310 80164
rect 55412 80052 55468 80108
rect 82012 80052 82068 80108
rect 55412 79996 69580 80052
rect 69636 79996 69646 80052
rect 82012 79996 85596 80052
rect 85652 79996 85820 80052
rect 85876 79996 85886 80052
rect 19826 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20110 79996
rect 50546 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50830 79996
rect 81266 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81550 79996
rect 88386 79884 88396 79940
rect 88452 79884 89628 79940
rect 89684 79884 95340 79940
rect 95396 79884 95406 79940
rect 52322 79772 52332 79828
rect 52388 79772 52892 79828
rect 52948 79772 55244 79828
rect 55300 79772 55310 79828
rect 56690 79772 56700 79828
rect 56756 79772 59500 79828
rect 59556 79772 59566 79828
rect 69570 79772 69580 79828
rect 69636 79772 72268 79828
rect 72324 79772 72334 79828
rect 86818 79772 86828 79828
rect 86884 79772 89180 79828
rect 89236 79772 89246 79828
rect 95666 79772 95676 79828
rect 95732 79772 97244 79828
rect 97300 79772 97310 79828
rect 54562 79660 54572 79716
rect 54628 79660 57372 79716
rect 57428 79660 57438 79716
rect 66434 79660 66444 79716
rect 66500 79660 70252 79716
rect 70308 79660 70318 79716
rect 80658 79660 80668 79716
rect 80724 79660 82124 79716
rect 82180 79660 82190 79716
rect 86258 79660 86268 79716
rect 86324 79660 87388 79716
rect 87444 79660 87454 79716
rect 91410 79660 91420 79716
rect 91476 79660 93772 79716
rect 93828 79660 94892 79716
rect 94948 79660 94958 79716
rect 95218 79660 95228 79716
rect 95284 79660 96124 79716
rect 96180 79660 96190 79716
rect 54674 79548 54684 79604
rect 54740 79548 55916 79604
rect 55972 79548 55982 79604
rect 56578 79548 56588 79604
rect 56644 79548 58268 79604
rect 58324 79548 58334 79604
rect 62626 79548 62636 79604
rect 62692 79548 63308 79604
rect 63364 79548 65660 79604
rect 65716 79548 65726 79604
rect 66780 79548 71484 79604
rect 71540 79548 71550 79604
rect 81442 79548 81452 79604
rect 81508 79548 83580 79604
rect 83636 79548 83646 79604
rect 84354 79548 84364 79604
rect 84420 79548 85484 79604
rect 85540 79548 86044 79604
rect 86100 79548 86110 79604
rect 96338 79548 96348 79604
rect 96404 79548 97580 79604
rect 97636 79548 97646 79604
rect 66780 79492 66836 79548
rect 57922 79436 57932 79492
rect 57988 79436 61180 79492
rect 61236 79436 66780 79492
rect 66836 79436 66846 79492
rect 77186 79436 77196 79492
rect 77252 79436 78876 79492
rect 78932 79436 78942 79492
rect 83122 79436 83132 79492
rect 83188 79436 84252 79492
rect 84308 79436 85260 79492
rect 85316 79436 85326 79492
rect 91858 79436 91868 79492
rect 91924 79436 92540 79492
rect 92596 79436 92606 79492
rect 56914 79324 56924 79380
rect 56980 79324 59500 79380
rect 59556 79324 59566 79380
rect 91634 79324 91644 79380
rect 91700 79324 93996 79380
rect 94052 79324 94062 79380
rect 83122 79212 83132 79268
rect 83188 79212 83468 79268
rect 83524 79212 83534 79268
rect 4466 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4750 79212
rect 35186 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35470 79212
rect 65906 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66190 79212
rect 96626 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96910 79212
rect 53666 78988 53676 79044
rect 53732 78988 54572 79044
rect 54628 78988 54638 79044
rect 59042 78988 59052 79044
rect 59108 78988 59118 79044
rect 78866 78988 78876 79044
rect 78932 78988 79884 79044
rect 79940 78988 80444 79044
rect 80500 78988 81788 79044
rect 81844 78988 81854 79044
rect 59052 78932 59108 78988
rect 58818 78876 58828 78932
rect 58884 78876 59108 78932
rect 66322 78876 66332 78932
rect 66388 78876 67228 78932
rect 67284 78876 67294 78932
rect 83570 78876 83580 78932
rect 83636 78876 87724 78932
rect 87780 78876 87790 78932
rect 90692 78876 94332 78932
rect 94388 78876 94398 78932
rect 90692 78820 90748 78876
rect 50194 78764 50204 78820
rect 50260 78764 52108 78820
rect 52164 78764 52174 78820
rect 53330 78764 53340 78820
rect 53396 78764 54236 78820
rect 54292 78764 54302 78820
rect 60386 78764 60396 78820
rect 60452 78764 62300 78820
rect 62356 78764 62366 78820
rect 66546 78764 66556 78820
rect 66612 78764 69804 78820
rect 69860 78764 69870 78820
rect 75180 78764 75740 78820
rect 75796 78764 75806 78820
rect 82786 78764 82796 78820
rect 82852 78764 84252 78820
rect 84308 78764 85932 78820
rect 85988 78764 85998 78820
rect 87490 78764 87500 78820
rect 87556 78764 90412 78820
rect 90468 78764 90748 78820
rect 75180 78708 75236 78764
rect 49298 78652 49308 78708
rect 49364 78652 50092 78708
rect 50148 78652 50764 78708
rect 50820 78652 50830 78708
rect 67778 78652 67788 78708
rect 67844 78652 69020 78708
rect 69076 78652 69086 78708
rect 71698 78652 71708 78708
rect 71764 78652 74172 78708
rect 74228 78652 75180 78708
rect 75236 78652 75246 78708
rect 75506 78652 75516 78708
rect 75572 78652 76300 78708
rect 76356 78652 76748 78708
rect 76804 78652 83356 78708
rect 83412 78652 83692 78708
rect 83748 78652 84140 78708
rect 84196 78652 84206 78708
rect 71708 78596 71764 78652
rect 49746 78540 49756 78596
rect 49812 78540 50204 78596
rect 50260 78540 50270 78596
rect 50978 78540 50988 78596
rect 51044 78540 52332 78596
rect 52388 78540 52398 78596
rect 57810 78540 57820 78596
rect 57876 78540 59724 78596
rect 59780 78540 61292 78596
rect 61348 78540 62972 78596
rect 63028 78540 63038 78596
rect 69346 78540 69356 78596
rect 69412 78540 70588 78596
rect 70644 78540 71764 78596
rect 88386 78540 88396 78596
rect 88452 78540 89516 78596
rect 89572 78540 95564 78596
rect 95620 78540 97804 78596
rect 97860 78540 97870 78596
rect 19826 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20110 78428
rect 50546 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50830 78428
rect 81266 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81550 78428
rect 58818 78316 58828 78372
rect 58884 78316 60956 78372
rect 61012 78316 61740 78372
rect 61796 78316 63420 78372
rect 63476 78316 67676 78372
rect 67732 78316 67742 78372
rect 48850 78204 48860 78260
rect 48916 78204 49644 78260
rect 49700 78204 49710 78260
rect 50418 78204 50428 78260
rect 50484 78204 67788 78260
rect 67844 78204 67854 78260
rect 68114 78204 68124 78260
rect 68180 78204 70028 78260
rect 70084 78204 70094 78260
rect 48290 78092 48300 78148
rect 48356 78092 49756 78148
rect 49812 78092 50316 78148
rect 50372 78092 51324 78148
rect 51380 78092 51390 78148
rect 76178 78092 76188 78148
rect 76244 78092 77308 78148
rect 77364 78092 77374 78148
rect 84578 78092 84588 78148
rect 84644 78092 89516 78148
rect 89572 78092 89582 78148
rect 50530 77980 50540 78036
rect 50596 77980 51772 78036
rect 51828 77980 52668 78036
rect 52724 77980 52734 78036
rect 58034 77980 58044 78036
rect 58100 77980 60060 78036
rect 60116 77980 60126 78036
rect 76738 77980 76748 78036
rect 76804 77980 78092 78036
rect 78148 77980 78158 78036
rect 87602 77980 87612 78036
rect 87668 77980 89180 78036
rect 89236 77980 89246 78036
rect 94434 77980 94444 78036
rect 94500 77980 95228 78036
rect 95284 77980 95294 78036
rect 51202 77868 51212 77924
rect 51268 77868 53116 77924
rect 53172 77868 53182 77924
rect 56690 77868 56700 77924
rect 56756 77868 57372 77924
rect 57428 77868 58156 77924
rect 58212 77868 58604 77924
rect 58660 77868 58670 77924
rect 72594 77868 72604 77924
rect 72660 77868 73164 77924
rect 73220 77868 73230 77924
rect 81330 77868 81340 77924
rect 81396 77868 82124 77924
rect 82180 77868 82190 77924
rect 72930 77756 72940 77812
rect 72996 77756 74956 77812
rect 75012 77756 75022 77812
rect 58370 77644 58380 77700
rect 58436 77644 61628 77700
rect 61684 77644 61694 77700
rect 4466 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4750 77644
rect 35186 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35470 77644
rect 65906 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66190 77644
rect 96626 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96910 77644
rect 68450 77420 68460 77476
rect 68516 77420 78540 77476
rect 78596 77420 78876 77476
rect 78932 77420 78942 77476
rect 50082 77308 50092 77364
rect 50148 77308 51996 77364
rect 52052 77308 52062 77364
rect 63074 77308 63084 77364
rect 63140 77308 70588 77364
rect 77746 77308 77756 77364
rect 77812 77308 79436 77364
rect 79492 77308 80780 77364
rect 80836 77308 80846 77364
rect 84354 77308 84364 77364
rect 84420 77308 85596 77364
rect 85652 77308 89404 77364
rect 89460 77308 89470 77364
rect 52322 77196 52332 77252
rect 52388 77196 52892 77252
rect 52948 77196 57708 77252
rect 57764 77196 62076 77252
rect 62132 77196 62972 77252
rect 63028 77196 67900 77252
rect 67956 77196 69580 77252
rect 69636 77196 69646 77252
rect 51650 77084 51660 77140
rect 51716 77084 54236 77140
rect 54292 77084 54302 77140
rect 70532 77028 70588 77308
rect 70802 77196 70812 77252
rect 70868 77196 71820 77252
rect 71876 77196 71886 77252
rect 73938 77196 73948 77252
rect 74004 77196 76524 77252
rect 76580 77196 76972 77252
rect 77028 77196 77038 77252
rect 78306 77196 78316 77252
rect 78372 77196 78988 77252
rect 79202 77196 79212 77252
rect 79268 77196 80444 77252
rect 80500 77196 84980 77252
rect 85250 77196 85260 77252
rect 85316 77196 86156 77252
rect 86212 77196 86222 77252
rect 78932 77140 78988 77196
rect 84924 77140 84980 77196
rect 72146 77084 72156 77140
rect 72212 77084 72716 77140
rect 72772 77084 72782 77140
rect 74722 77084 74732 77140
rect 74788 77084 77196 77140
rect 77252 77084 77262 77140
rect 78932 77084 82852 77140
rect 83010 77084 83020 77140
rect 83076 77084 84700 77140
rect 84756 77084 84766 77140
rect 84924 77084 86716 77140
rect 86772 77084 86782 77140
rect 49858 76972 49868 77028
rect 49924 76972 53340 77028
rect 53396 76972 53788 77028
rect 53844 76972 54348 77028
rect 54404 76972 54414 77028
rect 57362 76972 57372 77028
rect 57428 76972 58604 77028
rect 58660 76972 58670 77028
rect 58930 76972 58940 77028
rect 58996 76972 65436 77028
rect 65492 76972 66668 77028
rect 66724 76972 66734 77028
rect 70532 76972 72212 77028
rect 74274 76972 74284 77028
rect 74340 76972 75516 77028
rect 75572 76972 75582 77028
rect 78754 76972 78764 77028
rect 78820 76972 79212 77028
rect 79268 76972 79278 77028
rect 72156 76916 72212 76972
rect 82796 76916 82852 77084
rect 83346 76972 83356 77028
rect 83412 76972 84252 77028
rect 84308 76972 84318 77028
rect 94434 76972 94444 77028
rect 94500 76972 94780 77028
rect 94836 76972 95004 77028
rect 95060 76972 96012 77028
rect 96068 76972 97132 77028
rect 97188 76972 97198 77028
rect 72146 76860 72156 76916
rect 72212 76860 72222 76916
rect 82796 76860 85372 76916
rect 85428 76860 86044 76916
rect 86100 76860 86110 76916
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 81266 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81550 76860
rect 55234 76636 55244 76692
rect 55300 76636 58268 76692
rect 58324 76636 58334 76692
rect 63522 76636 63532 76692
rect 63588 76636 64540 76692
rect 64596 76636 67788 76692
rect 67844 76636 67854 76692
rect 75842 76636 75852 76692
rect 75908 76636 77756 76692
rect 77812 76636 78316 76692
rect 78372 76636 78382 76692
rect 80770 76636 80780 76692
rect 80836 76636 85708 76692
rect 85764 76636 85774 76692
rect 54226 76524 54236 76580
rect 54292 76524 54908 76580
rect 54964 76524 57596 76580
rect 57652 76524 58156 76580
rect 58212 76524 58222 76580
rect 64754 76524 64764 76580
rect 64820 76524 66444 76580
rect 66500 76524 66510 76580
rect 66658 76524 66668 76580
rect 66724 76524 67228 76580
rect 67284 76524 67294 76580
rect 75394 76524 75404 76580
rect 75460 76524 82796 76580
rect 82852 76524 82862 76580
rect 58482 76412 58492 76468
rect 58548 76412 58940 76468
rect 58996 76412 59006 76468
rect 66770 76412 66780 76468
rect 66836 76412 68124 76468
rect 68180 76412 70588 76468
rect 70644 76412 71260 76468
rect 71316 76412 71326 76468
rect 80546 76412 80556 76468
rect 80612 76412 82348 76468
rect 82404 76412 84308 76468
rect 84252 76356 84308 76412
rect 53778 76300 53788 76356
rect 53844 76300 56476 76356
rect 56532 76300 57372 76356
rect 57428 76300 57438 76356
rect 63858 76300 63868 76356
rect 63924 76300 64428 76356
rect 64484 76300 64494 76356
rect 71922 76300 71932 76356
rect 71988 76300 72604 76356
rect 72660 76300 74396 76356
rect 74452 76300 74462 76356
rect 84242 76300 84252 76356
rect 84308 76300 84318 76356
rect 85362 76300 85372 76356
rect 85428 76300 86380 76356
rect 86436 76300 86446 76356
rect 52658 76188 52668 76244
rect 52724 76188 53564 76244
rect 53620 76188 53630 76244
rect 66882 76188 66892 76244
rect 66948 76188 72828 76244
rect 72884 76188 73724 76244
rect 73780 76188 74284 76244
rect 74340 76188 74350 76244
rect 81554 76188 81564 76244
rect 81620 76188 82236 76244
rect 82292 76188 82302 76244
rect 72146 76076 72156 76132
rect 72212 76076 78764 76132
rect 78820 76076 78830 76132
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 96626 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96910 76076
rect 67218 75964 67228 76020
rect 67284 75964 67788 76020
rect 67844 75964 67854 76020
rect 61506 75852 61516 75908
rect 61572 75852 67340 75908
rect 67396 75852 67406 75908
rect 62962 75740 62972 75796
rect 63028 75740 63868 75796
rect 63924 75740 63934 75796
rect 64530 75740 64540 75796
rect 64596 75740 66444 75796
rect 66500 75740 66510 75796
rect 67172 75684 67228 75852
rect 71250 75740 71260 75796
rect 71316 75740 71596 75796
rect 71652 75740 71932 75796
rect 71988 75740 72044 75796
rect 72100 75740 72110 75796
rect 73378 75740 73388 75796
rect 73444 75740 74284 75796
rect 74340 75740 75404 75796
rect 75460 75740 75470 75796
rect 79762 75740 79772 75796
rect 79828 75740 81228 75796
rect 81284 75740 81294 75796
rect 86034 75740 86044 75796
rect 86100 75740 86716 75796
rect 86772 75740 86782 75796
rect 93538 75740 93548 75796
rect 93604 75740 95340 75796
rect 95396 75740 95406 75796
rect 66210 75628 66220 75684
rect 66276 75628 66892 75684
rect 66948 75628 66958 75684
rect 67172 75628 68012 75684
rect 68068 75628 71932 75684
rect 71988 75628 71998 75684
rect 73714 75628 73724 75684
rect 73780 75628 74788 75684
rect 74946 75628 74956 75684
rect 75012 75628 76300 75684
rect 76356 75628 77420 75684
rect 77476 75628 77486 75684
rect 81442 75628 81452 75684
rect 81508 75628 82348 75684
rect 82404 75628 82414 75684
rect 82786 75628 82796 75684
rect 82852 75628 83468 75684
rect 83524 75628 83534 75684
rect 84242 75628 84252 75684
rect 84308 75628 85260 75684
rect 85316 75628 85326 75684
rect 86370 75628 86380 75684
rect 86436 75628 86940 75684
rect 86996 75628 87006 75684
rect 94882 75628 94892 75684
rect 94948 75628 96012 75684
rect 96068 75628 96078 75684
rect 74732 75572 74788 75628
rect 74732 75516 75068 75572
rect 75124 75516 75134 75572
rect 75954 75516 75964 75572
rect 76020 75516 80556 75572
rect 80612 75516 80622 75572
rect 83234 75516 83244 75572
rect 83300 75516 84588 75572
rect 84644 75516 87052 75572
rect 87108 75516 87118 75572
rect 52658 75404 52668 75460
rect 52724 75404 55132 75460
rect 55188 75404 55198 75460
rect 82226 75404 82236 75460
rect 82292 75404 82572 75460
rect 82628 75404 84028 75460
rect 84084 75404 84094 75460
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 81266 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81550 75292
rect 51650 75180 51660 75236
rect 51716 75180 53340 75236
rect 53396 75180 54796 75236
rect 54852 75180 54862 75236
rect 90626 75180 90636 75236
rect 90692 75180 91420 75236
rect 91476 75180 91486 75236
rect 52210 75068 52220 75124
rect 52276 75068 54124 75124
rect 54180 75068 54190 75124
rect 54562 75068 54572 75124
rect 54628 75068 55692 75124
rect 55748 75068 55758 75124
rect 64418 75068 64428 75124
rect 64484 75068 65436 75124
rect 65492 75068 65502 75124
rect 69682 75068 69692 75124
rect 69748 75068 70588 75124
rect 70644 75068 70654 75124
rect 74610 75068 74620 75124
rect 74676 75068 75964 75124
rect 76020 75068 76030 75124
rect 78932 75068 98252 75124
rect 98308 75068 98318 75124
rect 78932 75012 78988 75068
rect 99200 75012 100000 75040
rect 50754 74956 50764 75012
rect 50820 74956 51884 75012
rect 51940 74956 51950 75012
rect 52882 74956 52892 75012
rect 52948 74956 54348 75012
rect 54404 74956 54414 75012
rect 74386 74956 74396 75012
rect 74452 74956 75068 75012
rect 75124 74956 78988 75012
rect 92306 74956 92316 75012
rect 92372 74956 93212 75012
rect 93268 74956 94332 75012
rect 94388 74956 94398 75012
rect 94546 74956 94556 75012
rect 94612 74956 100000 75012
rect 99200 74928 100000 74956
rect 54114 74844 54124 74900
rect 54180 74844 55916 74900
rect 55972 74844 55982 74900
rect 60610 74844 60620 74900
rect 60676 74844 64316 74900
rect 64372 74844 64382 74900
rect 73714 74844 73724 74900
rect 73780 74844 74284 74900
rect 74340 74844 74350 74900
rect 78418 74844 78428 74900
rect 78484 74844 84028 74900
rect 84084 74844 84094 74900
rect 88274 74844 88284 74900
rect 88340 74844 89404 74900
rect 89460 74844 89470 74900
rect 53666 74732 53676 74788
rect 53732 74732 54460 74788
rect 54516 74732 54796 74788
rect 54852 74732 55244 74788
rect 55300 74732 56476 74788
rect 56532 74732 61516 74788
rect 61572 74732 61582 74788
rect 89730 74732 89740 74788
rect 89796 74732 90860 74788
rect 90916 74732 92092 74788
rect 92148 74732 92158 74788
rect 93762 74732 93772 74788
rect 93828 74732 96348 74788
rect 96404 74732 96414 74788
rect 71698 74620 71708 74676
rect 71764 74620 72268 74676
rect 72324 74620 73500 74676
rect 73556 74620 89068 74676
rect 89124 74620 89964 74676
rect 90020 74620 90030 74676
rect 91746 74620 91756 74676
rect 91812 74620 92428 74676
rect 92484 74620 93548 74676
rect 93604 74620 93614 74676
rect 83010 74508 83020 74564
rect 83076 74508 83580 74564
rect 83636 74508 83646 74564
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 96626 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96910 74508
rect 91084 74284 91980 74340
rect 92036 74284 93100 74340
rect 93156 74284 93166 74340
rect 91084 74228 91140 74284
rect 50194 74172 50204 74228
rect 50260 74172 50652 74228
rect 50708 74172 52444 74228
rect 52500 74172 53116 74228
rect 53172 74172 53340 74228
rect 53396 74172 64428 74228
rect 64484 74172 64494 74228
rect 82226 74172 82236 74228
rect 82292 74172 82796 74228
rect 82852 74172 82862 74228
rect 89954 74172 89964 74228
rect 90020 74172 91084 74228
rect 91140 74172 91150 74228
rect 91634 74172 91644 74228
rect 91700 74172 92540 74228
rect 92596 74172 92606 74228
rect 96338 74172 96348 74228
rect 96404 74172 97804 74228
rect 97860 74172 97870 74228
rect 91644 74116 91700 74172
rect 60386 74060 60396 74116
rect 60452 74060 61516 74116
rect 61572 74060 61582 74116
rect 87826 74060 87836 74116
rect 87892 74060 89516 74116
rect 89572 74060 91700 74116
rect 57810 73948 57820 74004
rect 57876 73948 58156 74004
rect 58212 73948 59724 74004
rect 59780 73948 61852 74004
rect 61908 73948 61918 74004
rect 68562 73948 68572 74004
rect 68628 73948 69468 74004
rect 69524 73948 69534 74004
rect 70578 73948 70588 74004
rect 70644 73948 71484 74004
rect 71540 73948 71550 74004
rect 72258 73948 72268 74004
rect 72324 73948 72716 74004
rect 72772 73948 73276 74004
rect 73332 73948 73724 74004
rect 73780 73948 73790 74004
rect 89730 73948 89740 74004
rect 89796 73948 91308 74004
rect 91364 73948 91374 74004
rect 93986 73948 93996 74004
rect 94052 73948 95788 74004
rect 95844 73948 97132 74004
rect 97188 73948 97198 74004
rect 57138 73836 57148 73892
rect 57204 73836 58268 73892
rect 58324 73836 59500 73892
rect 59556 73836 70028 73892
rect 70084 73836 71260 73892
rect 71316 73836 71708 73892
rect 71764 73836 71774 73892
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 81266 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81550 73724
rect 61506 73500 61516 73556
rect 61572 73500 64092 73556
rect 64148 73500 65324 73556
rect 65380 73500 65548 73556
rect 65604 73500 67564 73556
rect 67620 73500 67630 73556
rect 78530 73500 78540 73556
rect 78596 73500 79324 73556
rect 79380 73500 79390 73556
rect 76514 73388 76524 73444
rect 76580 73388 77868 73444
rect 77924 73388 78764 73444
rect 78820 73388 93660 73444
rect 93716 73388 93996 73444
rect 94052 73388 94062 73444
rect 88498 73276 88508 73332
rect 88564 73276 89404 73332
rect 89460 73276 89470 73332
rect 91746 73276 91756 73332
rect 91812 73276 92316 73332
rect 92372 73276 92382 73332
rect 95218 73276 95228 73332
rect 95284 73276 97580 73332
rect 97636 73276 97646 73332
rect 51874 73164 51884 73220
rect 51940 73164 52332 73220
rect 52388 73164 53004 73220
rect 53060 73164 53070 73220
rect 56466 73164 56476 73220
rect 56532 73164 60844 73220
rect 60900 73164 62076 73220
rect 62132 73164 62142 73220
rect 69794 73164 69804 73220
rect 69860 73164 71148 73220
rect 71204 73164 71214 73220
rect 75954 73164 75964 73220
rect 76020 73164 77196 73220
rect 77252 73164 78316 73220
rect 78372 73164 78382 73220
rect 78978 73052 78988 73108
rect 79044 73052 79996 73108
rect 80052 73052 80062 73108
rect 62514 72940 62524 72996
rect 62580 72940 64764 72996
rect 64820 72940 64830 72996
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 96626 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96910 72940
rect 56354 72716 56364 72772
rect 56420 72716 58044 72772
rect 58100 72716 58110 72772
rect 53890 72492 53900 72548
rect 53956 72492 57820 72548
rect 57876 72492 58380 72548
rect 58436 72492 58446 72548
rect 60386 72492 60396 72548
rect 60452 72492 61740 72548
rect 61796 72492 61806 72548
rect 86594 72492 86604 72548
rect 86660 72492 87164 72548
rect 87220 72492 87230 72548
rect 94658 72492 94668 72548
rect 94724 72492 97692 72548
rect 97748 72492 97758 72548
rect 55458 72380 55468 72436
rect 55524 72380 56140 72436
rect 56196 72380 56206 72436
rect 70802 72380 70812 72436
rect 70868 72380 72156 72436
rect 72212 72380 72222 72436
rect 91746 72380 91756 72436
rect 91812 72380 94556 72436
rect 94612 72380 94622 72436
rect 54674 72268 54684 72324
rect 54740 72268 55244 72324
rect 55300 72268 56476 72324
rect 56532 72268 56542 72324
rect 64418 72268 64428 72324
rect 64484 72268 65436 72324
rect 65492 72268 65772 72324
rect 65828 72268 65838 72324
rect 75170 72268 75180 72324
rect 75236 72268 77196 72324
rect 77252 72268 79100 72324
rect 79156 72268 79166 72324
rect 83906 72268 83916 72324
rect 83972 72268 84476 72324
rect 84532 72268 84542 72324
rect 92530 72268 92540 72324
rect 92596 72268 94108 72324
rect 94164 72268 94174 72324
rect 62738 72156 62748 72212
rect 62804 72156 63644 72212
rect 63700 72156 63980 72212
rect 64036 72156 64204 72212
rect 64260 72156 65324 72212
rect 65380 72156 65390 72212
rect 74386 72156 74396 72212
rect 74452 72156 77420 72212
rect 77476 72156 78988 72212
rect 79044 72156 80332 72212
rect 80388 72156 81116 72212
rect 81172 72156 81182 72212
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 81266 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81550 72156
rect 72258 72044 72268 72100
rect 72324 72044 73836 72100
rect 73892 72044 73902 72100
rect 75618 72044 75628 72100
rect 75684 72044 76524 72100
rect 76580 72044 76590 72100
rect 49746 71932 49756 71988
rect 49812 71932 50428 71988
rect 50484 71932 50494 71988
rect 72594 71932 72604 71988
rect 72660 71932 73612 71988
rect 73668 71932 74844 71988
rect 74900 71932 74910 71988
rect 83010 71820 83020 71876
rect 83076 71820 85372 71876
rect 85428 71820 85438 71876
rect 89170 71708 89180 71764
rect 89236 71708 89852 71764
rect 89908 71708 90748 71764
rect 90692 71652 90748 71708
rect 51426 71596 51436 71652
rect 51492 71596 52108 71652
rect 52164 71596 52780 71652
rect 52836 71596 52846 71652
rect 56690 71596 56700 71652
rect 56756 71596 57260 71652
rect 57316 71596 58492 71652
rect 58548 71596 58558 71652
rect 62738 71596 62748 71652
rect 62804 71596 63196 71652
rect 63252 71596 63756 71652
rect 63812 71596 63822 71652
rect 65314 71596 65324 71652
rect 65380 71596 72044 71652
rect 72100 71596 73276 71652
rect 73332 71596 73342 71652
rect 73826 71596 73836 71652
rect 73892 71596 75068 71652
rect 75124 71596 76076 71652
rect 76132 71596 76636 71652
rect 76692 71596 76702 71652
rect 79986 71596 79996 71652
rect 80052 71596 80556 71652
rect 80612 71596 81564 71652
rect 81620 71596 81630 71652
rect 90692 71596 91868 71652
rect 91924 71596 95564 71652
rect 95620 71596 95630 71652
rect 50754 71484 50764 71540
rect 50820 71484 52556 71540
rect 52612 71484 52622 71540
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 96626 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96910 71372
rect 60946 71148 60956 71204
rect 61012 71148 74284 71204
rect 74340 71148 75628 71204
rect 75684 71148 75694 71204
rect 82338 71148 82348 71204
rect 82404 71148 84252 71204
rect 84308 71148 85708 71204
rect 85764 71148 85774 71204
rect 89282 71148 89292 71204
rect 89348 71148 90860 71204
rect 90916 71148 90926 71204
rect 91970 71148 91980 71204
rect 92036 71148 92988 71204
rect 93044 71148 93054 71204
rect 57922 71036 57932 71092
rect 57988 71036 59052 71092
rect 59108 71036 59500 71092
rect 59556 71036 59566 71092
rect 60610 71036 60620 71092
rect 60676 71036 62188 71092
rect 62244 71036 62254 71092
rect 62850 71036 62860 71092
rect 62916 71036 63308 71092
rect 63364 71036 64316 71092
rect 64372 71036 64382 71092
rect 68114 71036 68124 71092
rect 68180 71036 69580 71092
rect 69636 71036 71372 71092
rect 71428 71036 71438 71092
rect 90692 71036 91308 71092
rect 91364 71036 93660 71092
rect 93716 71036 95004 71092
rect 95060 71036 96460 71092
rect 96516 71036 96526 71092
rect 90692 70980 90748 71036
rect 73266 70924 73276 70980
rect 73332 70924 76076 70980
rect 76132 70924 88060 70980
rect 88116 70924 89404 70980
rect 89460 70924 90748 70980
rect 90850 70924 90860 70980
rect 90916 70924 91980 70980
rect 92036 70924 93100 70980
rect 93156 70924 93166 70980
rect 48178 70812 48188 70868
rect 48244 70812 49532 70868
rect 49588 70812 49598 70868
rect 68562 70812 68572 70868
rect 68628 70812 71484 70868
rect 71540 70812 71550 70868
rect 85652 70812 85932 70868
rect 85988 70812 85998 70868
rect 85652 70756 85708 70812
rect 48066 70700 48076 70756
rect 48132 70700 53340 70756
rect 53396 70700 53564 70756
rect 53620 70700 53630 70756
rect 66322 70700 66332 70756
rect 66388 70700 68236 70756
rect 68292 70700 68796 70756
rect 68852 70700 68862 70756
rect 81442 70700 81452 70756
rect 81508 70700 83020 70756
rect 83076 70700 84588 70756
rect 84644 70700 85708 70756
rect 57148 70588 57372 70644
rect 57428 70588 60284 70644
rect 60340 70588 60350 70644
rect 71362 70588 71372 70644
rect 71428 70588 72044 70644
rect 72100 70588 72110 70644
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 57148 70532 57204 70588
rect 81266 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81550 70588
rect 52098 70476 52108 70532
rect 52164 70476 52668 70532
rect 52724 70476 52734 70532
rect 53666 70476 53676 70532
rect 53732 70476 55132 70532
rect 55188 70476 56476 70532
rect 56532 70476 57204 70532
rect 67442 70476 67452 70532
rect 67508 70476 69132 70532
rect 69188 70476 69198 70532
rect 82898 70476 82908 70532
rect 82964 70476 83356 70532
rect 83412 70476 83692 70532
rect 83748 70476 83758 70532
rect 95452 70476 95676 70532
rect 95732 70476 95742 70532
rect 56242 70364 56252 70420
rect 56308 70364 58604 70420
rect 58660 70364 58670 70420
rect 60610 70364 60620 70420
rect 60676 70364 61516 70420
rect 61572 70364 62972 70420
rect 63028 70364 63868 70420
rect 63924 70364 64764 70420
rect 64820 70364 64830 70420
rect 95452 70308 95508 70476
rect 65314 70252 65324 70308
rect 65380 70252 66780 70308
rect 66836 70252 67788 70308
rect 67844 70252 67854 70308
rect 75506 70252 75516 70308
rect 75572 70252 76188 70308
rect 76244 70252 76254 70308
rect 95442 70252 95452 70308
rect 95508 70252 95518 70308
rect 52882 70140 52892 70196
rect 52948 70140 55580 70196
rect 55636 70140 58828 70196
rect 58884 70140 59276 70196
rect 59332 70140 60732 70196
rect 60788 70140 60798 70196
rect 81890 70140 81900 70196
rect 81956 70140 87164 70196
rect 87220 70140 89628 70196
rect 89684 70140 89694 70196
rect 96450 70140 96460 70196
rect 96516 70140 97692 70196
rect 97748 70140 97758 70196
rect 58706 70028 58716 70084
rect 58772 70028 59724 70084
rect 59780 70028 60956 70084
rect 61012 70028 61022 70084
rect 71026 70028 71036 70084
rect 71092 70028 72828 70084
rect 72884 70028 72894 70084
rect 77186 70028 77196 70084
rect 77252 70028 78316 70084
rect 78372 70028 78382 70084
rect 85362 70028 85372 70084
rect 85428 70028 85596 70084
rect 85652 70028 86268 70084
rect 86324 70028 87052 70084
rect 87108 70028 87118 70084
rect 95106 70028 95116 70084
rect 95172 70028 97132 70084
rect 97188 70028 97198 70084
rect 54562 69916 54572 69972
rect 54628 69916 57596 69972
rect 57652 69916 57662 69972
rect 89618 69916 89628 69972
rect 89684 69916 90972 69972
rect 91028 69916 91038 69972
rect 75170 69804 75180 69860
rect 75236 69804 75740 69860
rect 75796 69804 75806 69860
rect 86370 69804 86380 69860
rect 86436 69804 87164 69860
rect 87220 69804 87230 69860
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 96626 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96910 69804
rect 78642 69692 78652 69748
rect 78708 69692 85708 69748
rect 85764 69692 85774 69748
rect 56476 69580 57932 69636
rect 57988 69580 57998 69636
rect 68674 69580 68684 69636
rect 68740 69580 70252 69636
rect 70308 69580 70318 69636
rect 71474 69580 71484 69636
rect 71540 69580 72492 69636
rect 72548 69580 72558 69636
rect 56476 69524 56532 69580
rect 55682 69468 55692 69524
rect 55748 69468 56476 69524
rect 56532 69468 56542 69524
rect 57138 69468 57148 69524
rect 57204 69468 59836 69524
rect 59892 69468 60396 69524
rect 60452 69468 60462 69524
rect 67666 69468 67676 69524
rect 67732 69468 69244 69524
rect 69300 69468 69310 69524
rect 76262 69468 76300 69524
rect 76356 69468 76366 69524
rect 81218 69468 81228 69524
rect 81284 69468 81900 69524
rect 81956 69468 81966 69524
rect 84354 69468 84364 69524
rect 84420 69468 86044 69524
rect 86100 69468 86110 69524
rect 94882 69468 94892 69524
rect 94948 69468 95340 69524
rect 95396 69468 95676 69524
rect 95732 69468 95742 69524
rect 96002 69468 96012 69524
rect 96068 69468 97020 69524
rect 97076 69468 97086 69524
rect 48962 69356 48972 69412
rect 49028 69356 49532 69412
rect 49588 69356 52668 69412
rect 52724 69356 52734 69412
rect 65426 69356 65436 69412
rect 65492 69356 69356 69412
rect 69412 69356 69422 69412
rect 74946 69356 74956 69412
rect 75012 69356 75404 69412
rect 75460 69356 79100 69412
rect 79156 69356 79166 69412
rect 84466 69356 84476 69412
rect 84532 69356 89068 69412
rect 89124 69356 90300 69412
rect 90356 69356 90366 69412
rect 56466 69244 56476 69300
rect 56532 69244 57820 69300
rect 57876 69244 57886 69300
rect 71362 69244 71372 69300
rect 71428 69244 72380 69300
rect 72436 69244 73052 69300
rect 73108 69244 73118 69300
rect 74050 69244 74060 69300
rect 74116 69244 74844 69300
rect 74900 69244 77420 69300
rect 77476 69244 77486 69300
rect 78194 69244 78204 69300
rect 78260 69244 79996 69300
rect 80052 69244 80062 69300
rect 82114 69244 82124 69300
rect 82180 69244 82684 69300
rect 82740 69244 82750 69300
rect 88162 69244 88172 69300
rect 88228 69244 88844 69300
rect 88900 69244 88910 69300
rect 91634 69244 91644 69300
rect 91700 69244 93212 69300
rect 93268 69244 93278 69300
rect 52658 69132 52668 69188
rect 52724 69132 53676 69188
rect 53732 69132 53742 69188
rect 67330 69132 67340 69188
rect 67396 69132 68236 69188
rect 68292 69132 68302 69188
rect 76962 69132 76972 69188
rect 77028 69132 78540 69188
rect 78596 69132 78606 69188
rect 83570 69132 83580 69188
rect 83636 69132 84364 69188
rect 84420 69132 84430 69188
rect 74050 69020 74060 69076
rect 74116 69020 74732 69076
rect 74788 69020 74798 69076
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 81266 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81550 69020
rect 47842 68908 47852 68964
rect 47908 68908 50204 68964
rect 50260 68908 50270 68964
rect 60722 68908 60732 68964
rect 60788 68908 65436 68964
rect 65492 68908 65502 68964
rect 82562 68908 82572 68964
rect 82628 68908 83468 68964
rect 83524 68908 85260 68964
rect 85316 68908 85326 68964
rect 90514 68908 90524 68964
rect 90580 68908 93436 68964
rect 93492 68908 93502 68964
rect 51202 68796 51212 68852
rect 51268 68796 52780 68852
rect 52836 68796 53676 68852
rect 53732 68796 58716 68852
rect 58772 68796 58782 68852
rect 63634 68796 63644 68852
rect 63700 68796 70588 68852
rect 70644 68796 70654 68852
rect 74274 68796 74284 68852
rect 74340 68796 75180 68852
rect 75236 68796 75246 68852
rect 85810 68796 85820 68852
rect 85876 68796 87724 68852
rect 87780 68796 88732 68852
rect 88788 68796 88798 68852
rect 45938 68684 45948 68740
rect 46004 68684 54684 68740
rect 54740 68684 54750 68740
rect 73378 68684 73388 68740
rect 73444 68684 73500 68740
rect 73556 68684 73566 68740
rect 73714 68684 73724 68740
rect 73780 68684 75740 68740
rect 75796 68684 75806 68740
rect 78082 68684 78092 68740
rect 78148 68684 79100 68740
rect 79156 68684 79166 68740
rect 89506 68684 89516 68740
rect 89572 68684 90188 68740
rect 90244 68684 90254 68740
rect 49634 68572 49644 68628
rect 49700 68572 51884 68628
rect 51940 68572 51950 68628
rect 61506 68572 61516 68628
rect 61572 68572 62188 68628
rect 62244 68572 62254 68628
rect 63186 68572 63196 68628
rect 63252 68572 63532 68628
rect 63588 68572 63868 68628
rect 63924 68572 74284 68628
rect 74340 68572 74350 68628
rect 76290 68572 76300 68628
rect 76356 68572 77980 68628
rect 78036 68572 78046 68628
rect 83010 68572 83020 68628
rect 83076 68572 83916 68628
rect 83972 68572 87388 68628
rect 87444 68572 88508 68628
rect 88564 68572 91196 68628
rect 91252 68572 91868 68628
rect 91924 68572 91934 68628
rect 63196 68516 63252 68572
rect 62290 68460 62300 68516
rect 62356 68460 63252 68516
rect 67554 68460 67564 68516
rect 67620 68460 69916 68516
rect 69972 68460 71820 68516
rect 71876 68460 71886 68516
rect 50530 68348 50540 68404
rect 50596 68348 50988 68404
rect 51044 68348 53116 68404
rect 53172 68348 61852 68404
rect 61908 68348 62412 68404
rect 62468 68348 63196 68404
rect 63252 68348 63262 68404
rect 69570 68348 69580 68404
rect 69636 68348 74844 68404
rect 74900 68348 74910 68404
rect 79314 68348 79324 68404
rect 79380 68348 79996 68404
rect 80052 68348 80062 68404
rect 90178 68348 90188 68404
rect 90244 68348 92092 68404
rect 92148 68348 92158 68404
rect 67218 68236 67228 68292
rect 67284 68236 68348 68292
rect 68404 68236 68414 68292
rect 70578 68236 70588 68292
rect 70644 68236 72492 68292
rect 72548 68236 72558 68292
rect 73378 68236 73388 68292
rect 73444 68236 73724 68292
rect 73780 68236 73790 68292
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 96626 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96910 68236
rect 71334 68124 71372 68180
rect 71428 68124 73948 68180
rect 74004 68124 74014 68180
rect 62514 68012 62524 68068
rect 62580 68012 63420 68068
rect 63476 68012 63756 68068
rect 63812 68012 64316 68068
rect 64372 68012 64382 68068
rect 77970 68012 77980 68068
rect 78036 68012 90972 68068
rect 91028 68012 91038 68068
rect 75506 67900 75516 67956
rect 75572 67900 88956 67956
rect 89012 67900 89022 67956
rect 93538 67900 93548 67956
rect 93604 67900 95116 67956
rect 95172 67900 95182 67956
rect 66882 67788 66892 67844
rect 66948 67788 67452 67844
rect 67508 67788 67518 67844
rect 73826 67788 73836 67844
rect 73892 67732 73948 67844
rect 82562 67788 82572 67844
rect 82628 67788 83020 67844
rect 83076 67788 83086 67844
rect 83682 67788 83692 67844
rect 83748 67788 84252 67844
rect 84308 67788 84318 67844
rect 94658 67788 94668 67844
rect 94724 67788 96348 67844
rect 96404 67788 97356 67844
rect 97412 67788 98028 67844
rect 98084 67788 98094 67844
rect 60610 67676 60620 67732
rect 60676 67676 61516 67732
rect 61572 67676 61582 67732
rect 68450 67676 68460 67732
rect 68516 67676 69020 67732
rect 69076 67676 69086 67732
rect 73892 67676 74284 67732
rect 74340 67676 74350 67732
rect 75282 67676 75292 67732
rect 75348 67676 76300 67732
rect 76356 67676 77420 67732
rect 77476 67676 77486 67732
rect 85138 67676 85148 67732
rect 85204 67676 86044 67732
rect 86100 67676 86110 67732
rect 51090 67564 51100 67620
rect 51156 67564 52108 67620
rect 52164 67564 52174 67620
rect 52882 67564 52892 67620
rect 52948 67564 53340 67620
rect 53396 67564 53788 67620
rect 53844 67564 67564 67620
rect 67620 67564 67630 67620
rect 71558 67564 71596 67620
rect 71652 67564 71662 67620
rect 72034 67564 72044 67620
rect 72100 67564 72268 67620
rect 72324 67564 75068 67620
rect 75124 67564 75404 67620
rect 75460 67564 75470 67620
rect 79090 67564 79100 67620
rect 79156 67564 84308 67620
rect 85250 67564 85260 67620
rect 85316 67564 87500 67620
rect 87556 67564 87566 67620
rect 54226 67452 54236 67508
rect 54292 67452 68572 67508
rect 68628 67452 69580 67508
rect 69636 67452 69646 67508
rect 74470 67452 74508 67508
rect 74564 67452 74574 67508
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 81266 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81550 67452
rect 84252 67396 84308 67564
rect 68674 67340 68684 67396
rect 68740 67340 69916 67396
rect 69972 67340 69982 67396
rect 73350 67340 73388 67396
rect 73444 67340 73454 67396
rect 84242 67340 84252 67396
rect 84308 67340 84700 67396
rect 84756 67340 85820 67396
rect 85876 67340 85886 67396
rect 71596 67228 74508 67284
rect 74564 67228 75516 67284
rect 75572 67228 75582 67284
rect 83906 67228 83916 67284
rect 83972 67228 85372 67284
rect 85428 67228 85438 67284
rect 86482 67228 86492 67284
rect 86548 67228 88172 67284
rect 88228 67228 88238 67284
rect 71596 67172 71652 67228
rect 49746 67116 49756 67172
rect 49812 67116 51100 67172
rect 51156 67116 51884 67172
rect 51940 67116 53228 67172
rect 53284 67116 53788 67172
rect 53844 67116 53854 67172
rect 70242 67116 70252 67172
rect 70308 67116 70700 67172
rect 70756 67116 71652 67172
rect 73938 67116 73948 67172
rect 74004 67116 75740 67172
rect 75796 67116 75806 67172
rect 80098 67116 80108 67172
rect 80164 67116 81228 67172
rect 81284 67116 81294 67172
rect 82562 67116 82572 67172
rect 82628 67116 83244 67172
rect 83300 67116 83804 67172
rect 83860 67116 83870 67172
rect 85474 67116 85484 67172
rect 85540 67116 86716 67172
rect 86772 67116 87724 67172
rect 87780 67116 87790 67172
rect 88722 67116 88732 67172
rect 88788 67116 89068 67172
rect 89124 67116 89134 67172
rect 95442 67116 95452 67172
rect 95508 67116 96348 67172
rect 96404 67116 96414 67172
rect 48850 67004 48860 67060
rect 48916 67004 50428 67060
rect 50484 67004 52892 67060
rect 52948 67004 52958 67060
rect 77074 67004 77084 67060
rect 77140 67004 81564 67060
rect 81620 67004 83132 67060
rect 83188 67004 83580 67060
rect 83636 67004 83646 67060
rect 87826 67004 87836 67060
rect 87892 67004 90860 67060
rect 90916 67004 90926 67060
rect 91858 67004 91868 67060
rect 91924 67004 93996 67060
rect 94052 67004 95788 67060
rect 95844 67004 96908 67060
rect 96964 67004 96974 67060
rect 48290 66892 48300 66948
rect 48356 66892 49084 66948
rect 49140 66892 50204 66948
rect 50260 66892 50270 66948
rect 67442 66892 67452 66948
rect 67508 66892 69468 66948
rect 69524 66892 70140 66948
rect 70196 66892 70206 66948
rect 72146 66892 72156 66948
rect 72212 66892 73500 66948
rect 73556 66892 74732 66948
rect 74788 66892 75516 66948
rect 75572 66892 76748 66948
rect 76804 66892 76814 66948
rect 79202 66892 79212 66948
rect 79268 66892 80556 66948
rect 80612 66892 80622 66948
rect 93762 66892 93772 66948
rect 93828 66892 96012 66948
rect 96068 66892 97132 66948
rect 97188 66892 97198 66948
rect 54674 66780 54684 66836
rect 54740 66780 67788 66836
rect 67844 66780 67854 66836
rect 68786 66780 68796 66836
rect 68852 66780 71148 66836
rect 71204 66780 71214 66836
rect 80658 66780 80668 66836
rect 80724 66780 82012 66836
rect 82068 66780 82078 66836
rect 94098 66780 94108 66836
rect 94164 66780 95228 66836
rect 95284 66780 96124 66836
rect 96180 66780 97580 66836
rect 97636 66780 97646 66836
rect 71922 66668 71932 66724
rect 71988 66668 73948 66724
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 73892 66612 73948 66668
rect 96626 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96910 66668
rect 73892 66556 79100 66612
rect 79156 66556 79166 66612
rect 77410 66444 77420 66500
rect 77476 66444 81900 66500
rect 81956 66444 81966 66500
rect 82114 66444 82124 66500
rect 82180 66444 97468 66500
rect 97524 66444 97534 66500
rect 55234 66332 55244 66388
rect 55300 66332 56476 66388
rect 56532 66332 58044 66388
rect 58100 66332 58110 66388
rect 58268 66332 75964 66388
rect 76020 66332 76030 66388
rect 76188 66332 78652 66388
rect 78708 66332 78718 66388
rect 80770 66332 80780 66388
rect 80836 66332 82348 66388
rect 82404 66332 84028 66388
rect 84084 66332 84094 66388
rect 90962 66332 90972 66388
rect 91028 66332 94108 66388
rect 94164 66332 94174 66388
rect 58268 66276 58324 66332
rect 76188 66276 76244 66332
rect 52546 66220 52556 66276
rect 52612 66220 52892 66276
rect 52948 66220 52958 66276
rect 55794 66220 55804 66276
rect 55860 66220 58324 66276
rect 60386 66220 60396 66276
rect 60452 66220 61628 66276
rect 61684 66220 61694 66276
rect 66546 66220 66556 66276
rect 66612 66220 68572 66276
rect 68628 66220 68638 66276
rect 69794 66220 69804 66276
rect 69860 66220 73948 66276
rect 74050 66220 74060 66276
rect 74116 66220 76244 66276
rect 77634 66220 77644 66276
rect 77700 66220 78540 66276
rect 78596 66220 78606 66276
rect 85362 66220 85372 66276
rect 85428 66220 87052 66276
rect 87108 66220 87118 66276
rect 87378 66220 87388 66276
rect 87444 66220 87948 66276
rect 88004 66220 91532 66276
rect 91588 66220 91598 66276
rect 50194 66108 50204 66164
rect 50260 66108 51660 66164
rect 51716 66108 51726 66164
rect 58818 66108 58828 66164
rect 58884 66108 60508 66164
rect 60564 66108 60574 66164
rect 67890 66108 67900 66164
rect 67956 66108 69692 66164
rect 69748 66108 69758 66164
rect 70802 66108 70812 66164
rect 70868 66108 72492 66164
rect 72548 66108 73724 66164
rect 73780 66108 73790 66164
rect 73892 66052 73948 66220
rect 74732 66164 74788 66220
rect 74722 66108 74732 66164
rect 74788 66108 74798 66164
rect 74946 66108 74956 66164
rect 75012 66108 77756 66164
rect 77812 66108 77822 66164
rect 83234 66108 83244 66164
rect 83300 66108 84252 66164
rect 84308 66108 84318 66164
rect 90962 66108 90972 66164
rect 91028 66108 91420 66164
rect 91476 66108 91486 66164
rect 91308 66052 91364 66108
rect 49298 65996 49308 66052
rect 49364 65996 52220 66052
rect 52276 65996 52286 66052
rect 71026 65996 71036 66052
rect 71092 65996 72604 66052
rect 72660 65996 73276 66052
rect 73332 65996 73612 66052
rect 73668 65996 73678 66052
rect 73892 65996 77868 66052
rect 77924 65996 83580 66052
rect 83636 65996 84140 66052
rect 84196 65996 84206 66052
rect 85474 65996 85484 66052
rect 85540 65996 86492 66052
rect 86548 65996 87164 66052
rect 87220 65996 87230 66052
rect 90066 65996 90076 66052
rect 90132 65996 90860 66052
rect 90916 65996 90926 66052
rect 91298 65996 91308 66052
rect 91364 65996 91374 66052
rect 52322 65884 52332 65940
rect 52388 65884 54012 65940
rect 54068 65884 54078 65940
rect 62132 65884 69468 65940
rect 69524 65884 69804 65940
rect 69860 65884 69870 65940
rect 70924 65884 75740 65940
rect 75796 65884 75806 65940
rect 76178 65884 76188 65940
rect 76244 65884 77532 65940
rect 77588 65884 80668 65940
rect 80724 65884 80734 65940
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 62132 65828 62188 65884
rect 70924 65828 70980 65884
rect 81266 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81550 65884
rect 51762 65772 51772 65828
rect 51828 65772 52108 65828
rect 52164 65772 52444 65828
rect 52500 65772 52510 65828
rect 58818 65772 58828 65828
rect 58884 65772 59052 65828
rect 59108 65772 62188 65828
rect 66994 65772 67004 65828
rect 67060 65772 70924 65828
rect 70980 65772 70990 65828
rect 78530 65772 78540 65828
rect 78596 65772 81004 65828
rect 81060 65772 81070 65828
rect 82796 65772 85372 65828
rect 85428 65772 85438 65828
rect 88834 65772 88844 65828
rect 88900 65772 89068 65828
rect 89124 65772 90188 65828
rect 90244 65772 90254 65828
rect 82796 65716 82852 65772
rect 49186 65660 49196 65716
rect 49252 65660 50876 65716
rect 50932 65660 53340 65716
rect 53396 65660 53406 65716
rect 64978 65660 64988 65716
rect 65044 65660 65436 65716
rect 65492 65660 69244 65716
rect 69300 65660 69310 65716
rect 79090 65660 79100 65716
rect 79156 65660 80892 65716
rect 80948 65660 82796 65716
rect 82852 65660 82862 65716
rect 84354 65660 84364 65716
rect 84420 65660 86156 65716
rect 86212 65660 88060 65716
rect 88116 65660 88126 65716
rect 90300 65660 90860 65716
rect 90916 65660 90926 65716
rect 90300 65604 90356 65660
rect 50530 65548 50540 65604
rect 50596 65548 51436 65604
rect 51492 65548 51502 65604
rect 52434 65548 52444 65604
rect 52500 65548 53116 65604
rect 53172 65548 53182 65604
rect 54114 65548 54124 65604
rect 54180 65548 55020 65604
rect 55076 65548 55086 65604
rect 61842 65548 61852 65604
rect 61908 65548 62860 65604
rect 62916 65548 62926 65604
rect 64306 65548 64316 65604
rect 64372 65548 65660 65604
rect 65716 65548 65726 65604
rect 68908 65548 70700 65604
rect 70756 65548 70766 65604
rect 73042 65548 73052 65604
rect 73108 65548 73118 65604
rect 76066 65548 76076 65604
rect 76132 65548 79660 65604
rect 79716 65548 79726 65604
rect 80994 65548 81004 65604
rect 81060 65548 81900 65604
rect 81956 65548 81966 65604
rect 84130 65548 84140 65604
rect 84196 65548 86716 65604
rect 86772 65548 88284 65604
rect 88340 65548 88350 65604
rect 88946 65548 88956 65604
rect 89012 65548 89516 65604
rect 89572 65548 90300 65604
rect 90356 65548 90366 65604
rect 90626 65548 90636 65604
rect 90692 65548 91868 65604
rect 91924 65548 91934 65604
rect 96338 65548 96348 65604
rect 96404 65548 97580 65604
rect 97636 65548 97646 65604
rect 68908 65492 68964 65548
rect 73052 65492 73108 65548
rect 53676 65436 54572 65492
rect 54628 65436 55356 65492
rect 55412 65436 55804 65492
rect 55860 65436 55870 65492
rect 58930 65436 58940 65492
rect 58996 65436 59612 65492
rect 59668 65436 59678 65492
rect 66658 65436 66668 65492
rect 66724 65436 68964 65492
rect 71138 65436 71148 65492
rect 71204 65436 72604 65492
rect 72660 65436 72670 65492
rect 73052 65436 73948 65492
rect 74004 65436 74014 65492
rect 78418 65436 78428 65492
rect 78484 65436 79996 65492
rect 80052 65436 80062 65492
rect 88162 65436 88172 65492
rect 88228 65436 89180 65492
rect 89236 65436 89246 65492
rect 94322 65436 94332 65492
rect 94388 65436 95340 65492
rect 95396 65436 95406 65492
rect 53676 65268 53732 65436
rect 68338 65324 68348 65380
rect 68404 65324 72044 65380
rect 72100 65324 72110 65380
rect 72706 65324 72716 65380
rect 72772 65324 73724 65380
rect 73780 65324 73790 65380
rect 75394 65324 75404 65380
rect 75460 65324 78540 65380
rect 78596 65324 78606 65380
rect 80098 65324 80108 65380
rect 80164 65324 81116 65380
rect 81172 65324 81182 65380
rect 53666 65212 53676 65268
rect 53732 65212 53742 65268
rect 83010 65212 83020 65268
rect 83076 65212 86716 65268
rect 86772 65212 86782 65268
rect 67778 65100 67788 65156
rect 67844 65100 69692 65156
rect 69748 65100 79660 65156
rect 79716 65100 82236 65156
rect 82292 65100 82684 65156
rect 82740 65100 82796 65156
rect 82852 65100 82862 65156
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 96626 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96910 65100
rect 60834 64988 60844 65044
rect 60900 64988 62188 65044
rect 70354 64988 70364 65044
rect 70420 64988 78092 65044
rect 78148 64988 79436 65044
rect 79492 64988 80332 65044
rect 80388 64988 81228 65044
rect 81284 64988 81294 65044
rect 82870 64988 82908 65044
rect 82964 64988 82974 65044
rect 88498 64988 88508 65044
rect 88564 64988 93772 65044
rect 93828 64988 94220 65044
rect 94276 64988 95564 65044
rect 95620 64988 95630 65044
rect 62132 64932 62188 64988
rect 53442 64876 53452 64932
rect 53508 64876 54124 64932
rect 54180 64876 54190 64932
rect 62132 64876 67172 64932
rect 67330 64876 67340 64932
rect 67396 64876 68124 64932
rect 68180 64876 68460 64932
rect 68516 64876 70476 64932
rect 70532 64876 70542 64932
rect 70690 64876 70700 64932
rect 70756 64876 71260 64932
rect 71316 64876 72044 64932
rect 72100 64876 72110 64932
rect 78978 64876 78988 64932
rect 79044 64876 83580 64932
rect 83636 64876 83646 64932
rect 67116 64820 67172 64876
rect 27682 64764 27692 64820
rect 27748 64764 56364 64820
rect 56420 64764 56430 64820
rect 60498 64764 60508 64820
rect 60564 64764 61740 64820
rect 61796 64764 61806 64820
rect 62132 64764 67060 64820
rect 67116 64764 83132 64820
rect 83188 64764 83198 64820
rect 89394 64764 89404 64820
rect 89460 64764 90188 64820
rect 90244 64764 90748 64820
rect 90804 64764 90814 64820
rect 62132 64708 62188 64764
rect 67004 64708 67060 64764
rect 32162 64652 32172 64708
rect 32228 64652 46956 64708
rect 47012 64652 47022 64708
rect 50978 64652 50988 64708
rect 51044 64652 53340 64708
rect 53396 64652 53406 64708
rect 57586 64652 57596 64708
rect 57652 64652 58044 64708
rect 58100 64652 59500 64708
rect 59556 64652 59836 64708
rect 59892 64652 62188 64708
rect 64082 64652 64092 64708
rect 64148 64652 66332 64708
rect 66388 64652 66398 64708
rect 67004 64652 67340 64708
rect 67396 64652 67406 64708
rect 67666 64652 67676 64708
rect 67732 64652 71260 64708
rect 71316 64652 71326 64708
rect 71558 64652 71596 64708
rect 71652 64652 71662 64708
rect 74050 64652 74060 64708
rect 74116 64652 74396 64708
rect 74452 64652 74956 64708
rect 75012 64652 75022 64708
rect 79986 64652 79996 64708
rect 80052 64652 82684 64708
rect 82740 64652 83244 64708
rect 83300 64652 83310 64708
rect 97122 64652 97132 64708
rect 97188 64652 97692 64708
rect 97748 64652 97758 64708
rect 52434 64540 52444 64596
rect 52500 64540 53676 64596
rect 53732 64540 53742 64596
rect 54674 64540 54684 64596
rect 54740 64540 57484 64596
rect 57540 64540 57550 64596
rect 57810 64540 57820 64596
rect 57876 64540 59388 64596
rect 59444 64540 68236 64596
rect 68292 64540 68572 64596
rect 68628 64540 69356 64596
rect 69412 64540 69422 64596
rect 78306 64540 78316 64596
rect 78372 64540 78988 64596
rect 79044 64540 79054 64596
rect 80994 64540 81004 64596
rect 81060 64540 81788 64596
rect 81844 64540 88396 64596
rect 88452 64540 88462 64596
rect 56466 64428 56476 64484
rect 56532 64428 60284 64484
rect 60340 64428 60350 64484
rect 61730 64428 61740 64484
rect 61796 64428 73948 64484
rect 76850 64428 76860 64484
rect 76916 64428 77868 64484
rect 77924 64428 85484 64484
rect 85540 64428 85550 64484
rect 93650 64428 93660 64484
rect 93716 64428 94444 64484
rect 94500 64428 95564 64484
rect 95620 64428 95630 64484
rect 73892 64372 73948 64428
rect 55346 64316 55356 64372
rect 55412 64316 57596 64372
rect 57652 64316 58492 64372
rect 58548 64316 59276 64372
rect 59332 64316 61628 64372
rect 61684 64316 67340 64372
rect 67396 64316 67406 64372
rect 73892 64316 79324 64372
rect 79380 64316 79390 64372
rect 82786 64316 82796 64372
rect 82852 64316 88620 64372
rect 88676 64316 88686 64372
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 81266 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81550 64316
rect 56914 64204 56924 64260
rect 56980 64204 61964 64260
rect 62020 64204 62030 64260
rect 68898 64204 68908 64260
rect 68964 64204 79660 64260
rect 79716 64204 79884 64260
rect 79940 64204 79950 64260
rect 82450 64204 82460 64260
rect 82516 64204 85708 64260
rect 85652 64148 85708 64204
rect 57922 64092 57932 64148
rect 57988 64092 59052 64148
rect 59108 64092 59118 64148
rect 66210 64092 66220 64148
rect 66276 64092 71204 64148
rect 71698 64092 71708 64148
rect 71764 64092 72940 64148
rect 72996 64092 73006 64148
rect 77746 64092 77756 64148
rect 77812 64092 79100 64148
rect 79156 64092 79324 64148
rect 79380 64092 79390 64148
rect 79650 64092 79660 64148
rect 79716 64092 80220 64148
rect 80276 64092 80286 64148
rect 81106 64092 81116 64148
rect 81172 64092 82012 64148
rect 82068 64092 82078 64148
rect 82898 64092 82908 64148
rect 82964 64092 85540 64148
rect 85652 64092 86268 64148
rect 86324 64092 86334 64148
rect 86594 64092 86604 64148
rect 86660 64092 90300 64148
rect 90356 64092 90366 64148
rect 91298 64092 91308 64148
rect 91364 64092 93436 64148
rect 93492 64092 93502 64148
rect 94546 64092 94556 64148
rect 94612 64092 96348 64148
rect 96404 64092 96414 64148
rect 57474 63980 57484 64036
rect 57540 63980 58716 64036
rect 58772 63980 58940 64036
rect 58996 63980 59006 64036
rect 61180 63980 67004 64036
rect 67060 63980 67070 64036
rect 70578 63980 70588 64036
rect 70644 63980 70700 64036
rect 70756 63980 70766 64036
rect 61180 63924 61236 63980
rect 71148 63924 71204 64092
rect 85484 64036 85540 64092
rect 72034 63980 72044 64036
rect 72100 63980 72380 64036
rect 72436 63980 77084 64036
rect 77140 63980 77150 64036
rect 79986 63980 79996 64036
rect 80052 63980 81844 64036
rect 82786 63980 82796 64036
rect 82852 63980 84644 64036
rect 84802 63980 84812 64036
rect 84868 63980 85428 64036
rect 85484 63980 87612 64036
rect 87668 63980 87678 64036
rect 81788 63924 81844 63980
rect 84588 63924 84644 63980
rect 85372 63924 85428 63980
rect 52434 63868 52444 63924
rect 52500 63868 54236 63924
rect 54292 63868 54302 63924
rect 54460 63868 55020 63924
rect 55076 63868 55086 63924
rect 57922 63868 57932 63924
rect 57988 63868 61180 63924
rect 61236 63868 61246 63924
rect 61404 63868 66668 63924
rect 66724 63868 66734 63924
rect 67330 63868 67340 63924
rect 67396 63868 68348 63924
rect 68404 63868 68414 63924
rect 71148 63868 71708 63924
rect 71764 63868 71932 63924
rect 71988 63868 71998 63924
rect 72146 63868 72156 63924
rect 72212 63868 72716 63924
rect 72772 63868 72782 63924
rect 72930 63868 72940 63924
rect 72996 63868 74956 63924
rect 75012 63868 75404 63924
rect 75460 63868 75470 63924
rect 76402 63868 76412 63924
rect 76468 63868 77196 63924
rect 77252 63868 77980 63924
rect 78036 63868 78046 63924
rect 80434 63868 80444 63924
rect 80500 63868 81564 63924
rect 81620 63868 81630 63924
rect 81778 63868 81788 63924
rect 81844 63868 81854 63924
rect 82124 63868 82796 63924
rect 82852 63868 82862 63924
rect 83132 63868 83580 63924
rect 83636 63868 83916 63924
rect 83972 63868 83982 63924
rect 84588 63868 84924 63924
rect 84980 63868 84990 63924
rect 85138 63868 85148 63924
rect 85204 63868 85214 63924
rect 85372 63868 85932 63924
rect 85988 63868 85998 63924
rect 86258 63868 86268 63924
rect 86324 63868 87388 63924
rect 87444 63868 87454 63924
rect 89282 63868 89292 63924
rect 89348 63868 90412 63924
rect 90468 63868 92988 63924
rect 93044 63868 93054 63924
rect 54460 63812 54516 63868
rect 61404 63812 61460 63868
rect 48850 63756 48860 63812
rect 48916 63756 49532 63812
rect 49588 63756 49598 63812
rect 53442 63756 53452 63812
rect 53508 63756 54516 63812
rect 60386 63756 60396 63812
rect 60452 63756 61460 63812
rect 72258 63756 72268 63812
rect 72324 63756 72604 63812
rect 72660 63756 75964 63812
rect 76020 63756 76030 63812
rect 78754 63756 78764 63812
rect 78820 63756 79884 63812
rect 79940 63756 79950 63812
rect 82124 63700 82180 63868
rect 82870 63756 82908 63812
rect 82964 63756 82974 63812
rect 83132 63700 83188 63868
rect 85148 63700 85204 63868
rect 85362 63756 85372 63812
rect 85428 63756 86044 63812
rect 86100 63756 86110 63812
rect 90850 63756 90860 63812
rect 90916 63756 92540 63812
rect 92596 63756 92606 63812
rect 12562 63644 12572 63700
rect 12628 63644 62188 63700
rect 70690 63644 70700 63700
rect 70756 63644 70766 63700
rect 70914 63644 70924 63700
rect 70980 63644 71372 63700
rect 71428 63644 71438 63700
rect 75170 63644 75180 63700
rect 75236 63644 75460 63700
rect 75730 63644 75740 63700
rect 75796 63644 77868 63700
rect 77924 63644 77934 63700
rect 79650 63644 79660 63700
rect 79716 63644 82180 63700
rect 82758 63644 82796 63700
rect 82852 63644 82862 63700
rect 83122 63644 83132 63700
rect 83188 63644 83198 63700
rect 85148 63644 87052 63700
rect 87108 63644 87118 63700
rect 89506 63644 89516 63700
rect 89572 63644 90748 63700
rect 90804 63644 91196 63700
rect 91252 63644 91262 63700
rect 46946 63532 46956 63588
rect 47012 63532 59500 63588
rect 59556 63532 59566 63588
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 50306 63420 50316 63476
rect 50372 63420 52780 63476
rect 52836 63420 52846 63476
rect 52994 63420 53004 63476
rect 53060 63420 55692 63476
rect 55748 63420 55758 63476
rect 56354 63420 56364 63476
rect 56420 63420 57596 63476
rect 57652 63420 57662 63476
rect 62132 63364 62188 63644
rect 70700 63588 70756 63644
rect 75404 63588 75460 63644
rect 70700 63532 71036 63588
rect 71092 63532 71102 63588
rect 75394 63532 75404 63588
rect 75460 63532 75470 63588
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 96626 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96910 63532
rect 75506 63420 75516 63476
rect 75572 63420 76524 63476
rect 76580 63420 76590 63476
rect 50372 63308 54292 63364
rect 54450 63308 54460 63364
rect 54516 63308 57372 63364
rect 57428 63308 57438 63364
rect 57698 63308 57708 63364
rect 57764 63308 58156 63364
rect 58212 63308 58222 63364
rect 62132 63308 66220 63364
rect 66276 63308 66556 63364
rect 66612 63308 66622 63364
rect 76066 63308 76076 63364
rect 76132 63308 77756 63364
rect 77812 63308 77822 63364
rect 79314 63308 79324 63364
rect 79380 63308 82348 63364
rect 82404 63308 82414 63364
rect 88386 63308 88396 63364
rect 88452 63308 88956 63364
rect 89012 63308 89516 63364
rect 89572 63308 89582 63364
rect 50372 63252 50428 63308
rect 54236 63252 54292 63308
rect 47954 63196 47964 63252
rect 48020 63196 50428 63252
rect 52658 63196 52668 63252
rect 52724 63196 53340 63252
rect 53396 63196 53406 63252
rect 54236 63196 58268 63252
rect 58324 63196 58334 63252
rect 75954 63196 75964 63252
rect 76020 63196 77308 63252
rect 77364 63196 77374 63252
rect 79202 63196 79212 63252
rect 79268 63196 80668 63252
rect 80724 63196 80734 63252
rect 81554 63196 81564 63252
rect 81620 63196 84364 63252
rect 84420 63196 84430 63252
rect 86146 63196 86156 63252
rect 86212 63196 88732 63252
rect 88788 63196 88798 63252
rect 90066 63196 90076 63252
rect 90132 63196 92204 63252
rect 92260 63196 92270 63252
rect 52210 63084 52220 63140
rect 52276 63084 53564 63140
rect 53620 63084 54460 63140
rect 54516 63084 54526 63140
rect 56914 63084 56924 63140
rect 56980 63084 58940 63140
rect 58996 63084 59006 63140
rect 78530 63084 78540 63140
rect 78596 63084 83020 63140
rect 83076 63084 83086 63140
rect 85250 63084 85260 63140
rect 85316 63084 86268 63140
rect 86324 63084 86334 63140
rect 88386 63084 88396 63140
rect 88452 63084 89628 63140
rect 89684 63084 89694 63140
rect 91186 63084 91196 63140
rect 91252 63084 95004 63140
rect 95060 63084 96460 63140
rect 96516 63084 96526 63140
rect 31892 62972 69244 63028
rect 69300 62972 69916 63028
rect 69972 62972 69982 63028
rect 78754 62972 78764 63028
rect 78820 62972 81004 63028
rect 81060 62972 81070 63028
rect 83020 62972 83804 63028
rect 83860 62972 83870 63028
rect 84466 62972 84476 63028
rect 84532 62972 86044 63028
rect 86100 62972 86110 63028
rect 86594 62972 86604 63028
rect 86660 62972 90300 63028
rect 90356 62972 90366 63028
rect 31892 62916 31948 62972
rect 83020 62916 83076 62972
rect 8372 62860 31948 62916
rect 49410 62860 49420 62916
rect 49476 62860 51772 62916
rect 51828 62860 51838 62916
rect 58818 62860 58828 62916
rect 58884 62860 62188 62916
rect 62244 62860 62254 62916
rect 65874 62860 65884 62916
rect 65940 62860 66892 62916
rect 66948 62860 67116 62916
rect 67172 62860 67182 62916
rect 76514 62860 76524 62916
rect 76580 62860 79548 62916
rect 79604 62860 79614 62916
rect 80658 62860 80668 62916
rect 80724 62860 83020 62916
rect 83076 62860 83086 62916
rect 8372 62804 8428 62860
rect 83692 62804 83748 62972
rect 83906 62860 83916 62916
rect 83972 62860 85820 62916
rect 85876 62860 85886 62916
rect 88050 62860 88060 62916
rect 88116 62860 91756 62916
rect 91812 62860 91822 62916
rect 92306 62860 92316 62916
rect 92372 62860 94220 62916
rect 94276 62860 97020 62916
rect 97076 62860 97086 62916
rect 2146 62748 2156 62804
rect 2212 62748 8428 62804
rect 59266 62748 59276 62804
rect 59332 62748 60284 62804
rect 60340 62748 68908 62804
rect 68964 62748 68974 62804
rect 74386 62748 74396 62804
rect 74452 62748 74732 62804
rect 74788 62748 74798 62804
rect 83692 62748 86940 62804
rect 86996 62748 87006 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 81266 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81550 62748
rect 54114 62636 54124 62692
rect 54180 62636 56700 62692
rect 56756 62636 57036 62692
rect 57092 62636 71036 62692
rect 71092 62636 71932 62692
rect 71988 62636 75852 62692
rect 75908 62636 75918 62692
rect 82226 62636 82236 62692
rect 82292 62636 82684 62692
rect 82740 62636 82750 62692
rect 83020 62636 85148 62692
rect 85204 62636 87276 62692
rect 87332 62636 87948 62692
rect 88004 62636 88014 62692
rect 88162 62636 88172 62692
rect 88228 62636 93660 62692
rect 93716 62636 94332 62692
rect 94388 62636 95116 62692
rect 95172 62636 95676 62692
rect 95732 62636 97244 62692
rect 97300 62636 97310 62692
rect 83020 62580 83076 62636
rect 55122 62524 55132 62580
rect 55188 62524 58604 62580
rect 58660 62524 58670 62580
rect 60050 62524 60060 62580
rect 60116 62524 63308 62580
rect 63364 62524 63374 62580
rect 63970 62524 63980 62580
rect 64036 62524 76860 62580
rect 76916 62524 76926 62580
rect 80546 62524 80556 62580
rect 80612 62524 81900 62580
rect 81956 62524 83076 62580
rect 83234 62524 83244 62580
rect 83300 62524 84364 62580
rect 84420 62524 84430 62580
rect 84690 62524 84700 62580
rect 84756 62524 86828 62580
rect 86884 62524 86894 62580
rect 0 62468 800 62496
rect 63980 62468 64036 62524
rect 0 62412 1820 62468
rect 1876 62412 1886 62468
rect 51762 62412 51772 62468
rect 51828 62412 52668 62468
rect 52724 62412 52734 62468
rect 62178 62412 62188 62468
rect 62244 62412 63196 62468
rect 63252 62412 63420 62468
rect 63476 62412 64036 62468
rect 74498 62412 74508 62468
rect 74564 62412 74844 62468
rect 74900 62412 74910 62468
rect 79090 62412 79100 62468
rect 79156 62412 79436 62468
rect 79492 62412 79502 62468
rect 80322 62412 80332 62468
rect 80388 62412 81340 62468
rect 81396 62412 81406 62468
rect 81676 62412 82460 62468
rect 82516 62412 82526 62468
rect 83542 62412 83580 62468
rect 83636 62412 83646 62468
rect 84018 62412 84028 62468
rect 84084 62412 86548 62468
rect 87826 62412 87836 62468
rect 87892 62412 89068 62468
rect 89124 62412 89134 62468
rect 89282 62412 89292 62468
rect 89348 62412 93100 62468
rect 93156 62412 93166 62468
rect 0 62384 800 62412
rect 81676 62356 81732 62412
rect 86492 62356 86548 62412
rect 57810 62300 57820 62356
rect 57876 62300 58604 62356
rect 58660 62300 58670 62356
rect 70130 62300 70140 62356
rect 70196 62300 70476 62356
rect 70532 62300 71036 62356
rect 71092 62300 74508 62356
rect 74564 62300 75404 62356
rect 75460 62300 75628 62356
rect 75684 62300 75694 62356
rect 81666 62300 81676 62356
rect 81732 62300 81742 62356
rect 82114 62300 82124 62356
rect 82180 62300 83244 62356
rect 83300 62300 83310 62356
rect 83654 62300 83692 62356
rect 83748 62300 83758 62356
rect 83906 62300 83916 62356
rect 83972 62300 86044 62356
rect 86100 62300 86110 62356
rect 86482 62300 86492 62356
rect 86548 62300 86558 62356
rect 88610 62300 88620 62356
rect 88676 62300 89516 62356
rect 89572 62300 89582 62356
rect 92306 62300 92316 62356
rect 92372 62300 96348 62356
rect 96404 62300 96414 62356
rect 48850 62188 48860 62244
rect 48916 62188 50316 62244
rect 50372 62188 50382 62244
rect 64866 62188 64876 62244
rect 64932 62188 65772 62244
rect 65828 62188 65838 62244
rect 69906 62188 69916 62244
rect 69972 62188 70924 62244
rect 70980 62188 70990 62244
rect 71362 62188 71372 62244
rect 71428 62188 71484 62244
rect 71540 62188 74060 62244
rect 74116 62188 74126 62244
rect 79762 62188 79772 62244
rect 79828 62188 80780 62244
rect 80836 62188 83300 62244
rect 83458 62188 83468 62244
rect 83524 62188 85708 62244
rect 85764 62188 85774 62244
rect 91522 62188 91532 62244
rect 91588 62188 93212 62244
rect 93268 62188 93278 62244
rect 83244 62132 83300 62188
rect 71138 62076 71148 62132
rect 71204 62076 71708 62132
rect 71764 62076 75404 62132
rect 75460 62076 75470 62132
rect 75730 62076 75740 62132
rect 75796 62076 78092 62132
rect 78148 62076 78158 62132
rect 81666 62076 81676 62132
rect 81732 62076 82796 62132
rect 82852 62076 82862 62132
rect 83244 62076 83580 62132
rect 83636 62076 83646 62132
rect 72482 61964 72492 62020
rect 72548 61964 74396 62020
rect 74452 61964 78876 62020
rect 78932 61964 78942 62020
rect 79650 61964 79660 62020
rect 79716 61964 80108 62020
rect 80164 61964 80174 62020
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 96626 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96910 61964
rect 61842 61852 61852 61908
rect 61908 61852 62860 61908
rect 62916 61852 62926 61908
rect 72370 61852 72380 61908
rect 72436 61852 72828 61908
rect 72884 61852 72894 61908
rect 73266 61852 73276 61908
rect 73332 61852 74284 61908
rect 74340 61852 76300 61908
rect 76356 61852 80220 61908
rect 80276 61852 80286 61908
rect 69234 61740 69244 61796
rect 69300 61740 81452 61796
rect 81508 61740 86268 61796
rect 86324 61740 86334 61796
rect 83692 61684 83748 61740
rect 62738 61628 62748 61684
rect 62804 61628 63756 61684
rect 63812 61628 65996 61684
rect 66052 61628 66062 61684
rect 66546 61628 66556 61684
rect 66612 61628 68236 61684
rect 68292 61628 68460 61684
rect 68516 61628 68526 61684
rect 75394 61628 75404 61684
rect 75460 61628 82236 61684
rect 82292 61628 82302 61684
rect 83682 61628 83692 61684
rect 83748 61628 83758 61684
rect 85474 61628 85484 61684
rect 85540 61628 87612 61684
rect 87668 61628 87678 61684
rect 93202 61628 93212 61684
rect 93268 61628 95452 61684
rect 95508 61628 95518 61684
rect 55412 61516 56140 61572
rect 56196 61516 56206 61572
rect 62962 61516 62972 61572
rect 63028 61516 67452 61572
rect 67508 61516 69692 61572
rect 69748 61516 69758 61572
rect 70242 61516 70252 61572
rect 70308 61516 71148 61572
rect 71204 61516 72268 61572
rect 72324 61516 72334 61572
rect 75618 61516 75628 61572
rect 75684 61516 77308 61572
rect 77364 61516 77374 61572
rect 83458 61516 83468 61572
rect 83524 61516 83580 61572
rect 83636 61516 85260 61572
rect 85316 61516 85326 61572
rect 85652 61516 88284 61572
rect 88340 61516 89628 61572
rect 89684 61516 89694 61572
rect 55412 61460 55468 61516
rect 85652 61460 85708 61516
rect 55010 61404 55020 61460
rect 55076 61404 55468 61460
rect 55682 61404 55692 61460
rect 55748 61404 59164 61460
rect 59220 61404 60172 61460
rect 60228 61404 67676 61460
rect 67732 61404 69244 61460
rect 69300 61404 69310 61460
rect 70466 61404 70476 61460
rect 70532 61404 72828 61460
rect 72884 61404 76972 61460
rect 77028 61404 77038 61460
rect 77970 61404 77980 61460
rect 78036 61404 78988 61460
rect 79044 61404 85708 61460
rect 92530 61404 92540 61460
rect 92596 61404 94668 61460
rect 94724 61404 94734 61460
rect 55692 61348 55748 61404
rect 52322 61292 52332 61348
rect 52388 61292 53340 61348
rect 53396 61292 53406 61348
rect 55122 61292 55132 61348
rect 55188 61292 55748 61348
rect 56130 61292 56140 61348
rect 56196 61292 57036 61348
rect 57092 61292 57102 61348
rect 59266 61292 59276 61348
rect 59332 61292 59724 61348
rect 59780 61292 61628 61348
rect 61684 61292 61694 61348
rect 75170 61292 75180 61348
rect 75236 61292 77420 61348
rect 77476 61292 77486 61348
rect 79426 61292 79436 61348
rect 79492 61292 79502 61348
rect 79622 61292 79660 61348
rect 79716 61292 79726 61348
rect 81116 61292 84364 61348
rect 84420 61292 84430 61348
rect 84578 61292 84588 61348
rect 84644 61292 87164 61348
rect 87220 61292 87230 61348
rect 79436 61236 79492 61292
rect 81116 61236 81172 61292
rect 70018 61180 70028 61236
rect 70084 61180 70700 61236
rect 70756 61180 70766 61236
rect 72930 61180 72940 61236
rect 72996 61180 76300 61236
rect 76356 61180 76366 61236
rect 79436 61180 81172 61236
rect 91858 61180 91868 61236
rect 91924 61180 93324 61236
rect 93380 61180 93390 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 81266 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81550 61180
rect 59714 61068 59724 61124
rect 59780 61068 60396 61124
rect 60452 61068 60462 61124
rect 63634 61068 63644 61124
rect 63700 61068 66220 61124
rect 66276 61068 66286 61124
rect 84242 61068 84252 61124
rect 84308 61068 85820 61124
rect 85876 61068 85886 61124
rect 64082 60956 64092 61012
rect 64148 60956 66668 61012
rect 66724 60956 66734 61012
rect 77858 60956 77868 61012
rect 77924 60956 78876 61012
rect 78932 60956 79660 61012
rect 79716 60956 82404 61012
rect 82348 60900 82404 60956
rect 83244 60956 91644 61012
rect 91700 60956 91710 61012
rect 48402 60844 48412 60900
rect 48468 60844 49420 60900
rect 49476 60844 49486 60900
rect 61842 60844 61852 60900
rect 61908 60844 62300 60900
rect 62356 60844 65324 60900
rect 65380 60844 65548 60900
rect 65604 60844 69916 60900
rect 69972 60844 69982 60900
rect 70130 60844 70140 60900
rect 70196 60844 71372 60900
rect 71428 60844 72156 60900
rect 72212 60844 72492 60900
rect 72548 60844 72558 60900
rect 79314 60844 79324 60900
rect 79380 60844 81676 60900
rect 81732 60844 81742 60900
rect 82338 60844 82348 60900
rect 82404 60844 82796 60900
rect 82852 60844 82862 60900
rect 83244 60788 83300 60956
rect 84130 60844 84140 60900
rect 84196 60844 84588 60900
rect 84644 60844 84654 60900
rect 91644 60844 92428 60900
rect 92484 60844 92494 60900
rect 50418 60732 50428 60788
rect 50484 60732 50764 60788
rect 50820 60732 51100 60788
rect 51156 60732 51884 60788
rect 51940 60732 51950 60788
rect 56130 60732 56140 60788
rect 56196 60732 57372 60788
rect 57428 60732 57438 60788
rect 64530 60732 64540 60788
rect 64596 60732 65884 60788
rect 65940 60732 65950 60788
rect 67106 60732 67116 60788
rect 67172 60732 67676 60788
rect 67732 60732 67742 60788
rect 69346 60732 69356 60788
rect 69412 60732 70028 60788
rect 70084 60732 73500 60788
rect 73556 60732 73566 60788
rect 78754 60732 78764 60788
rect 78820 60732 83244 60788
rect 83300 60732 83310 60788
rect 84242 60732 84252 60788
rect 84308 60732 85708 60788
rect 85764 60732 85774 60788
rect 87042 60732 87052 60788
rect 87108 60732 89740 60788
rect 89796 60732 90748 60788
rect 90692 60676 90748 60732
rect 91644 60676 91700 60844
rect 50866 60620 50876 60676
rect 50932 60620 51436 60676
rect 51492 60620 52444 60676
rect 52500 60620 52510 60676
rect 60386 60620 60396 60676
rect 60452 60620 63980 60676
rect 64036 60620 76748 60676
rect 76804 60620 85596 60676
rect 85652 60620 86604 60676
rect 86660 60620 86670 60676
rect 86828 60620 88508 60676
rect 88564 60620 88574 60676
rect 90692 60620 91700 60676
rect 91756 60732 98140 60788
rect 98196 60732 98206 60788
rect 86828 60564 86884 60620
rect 91756 60564 91812 60732
rect 47618 60508 47628 60564
rect 47684 60508 49756 60564
rect 49812 60508 49822 60564
rect 63522 60508 63532 60564
rect 63588 60508 64876 60564
rect 64932 60508 64942 60564
rect 68002 60508 68012 60564
rect 68068 60508 69244 60564
rect 69300 60508 69310 60564
rect 70690 60508 70700 60564
rect 70756 60508 71484 60564
rect 71540 60508 71550 60564
rect 72146 60508 72156 60564
rect 72212 60508 73276 60564
rect 73332 60508 73342 60564
rect 73836 60508 80220 60564
rect 80276 60508 82236 60564
rect 82292 60508 82302 60564
rect 85586 60508 85596 60564
rect 85652 60508 86884 60564
rect 87938 60508 87948 60564
rect 88004 60508 89292 60564
rect 89348 60508 91812 60564
rect 92194 60508 92204 60564
rect 92260 60508 94108 60564
rect 94164 60508 94174 60564
rect 73836 60452 73892 60508
rect 67554 60396 67564 60452
rect 67620 60396 68460 60452
rect 68516 60396 69804 60452
rect 69860 60396 73892 60452
rect 75282 60396 75292 60452
rect 75348 60396 77532 60452
rect 77588 60396 79996 60452
rect 80052 60396 81452 60452
rect 81508 60396 81518 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 96626 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96910 60396
rect 72258 60284 72268 60340
rect 72324 60284 72716 60340
rect 72772 60284 72782 60340
rect 79650 60284 79660 60340
rect 79716 60284 83580 60340
rect 83636 60284 84028 60340
rect 84084 60284 84094 60340
rect 55570 60172 55580 60228
rect 55636 60172 57260 60228
rect 57316 60172 57326 60228
rect 71922 60172 71932 60228
rect 71988 60172 72940 60228
rect 72996 60172 73006 60228
rect 76962 60172 76972 60228
rect 77028 60172 77644 60228
rect 77700 60172 81340 60228
rect 81396 60172 83916 60228
rect 83972 60172 83982 60228
rect 50082 60060 50092 60116
rect 50148 60060 51212 60116
rect 51268 60060 51278 60116
rect 63634 60060 63644 60116
rect 63700 60060 67228 60116
rect 67284 60060 67294 60116
rect 69906 60060 69916 60116
rect 69972 60060 75852 60116
rect 75908 60060 76524 60116
rect 76580 60060 76590 60116
rect 79762 60060 79772 60116
rect 79828 60060 83132 60116
rect 83188 60060 85148 60116
rect 85204 60060 85214 60116
rect 48402 59948 48412 60004
rect 48468 59948 51772 60004
rect 51828 59948 52780 60004
rect 52836 59948 53676 60004
rect 53732 59948 53742 60004
rect 63074 59948 63084 60004
rect 63140 59948 64428 60004
rect 64484 59948 67340 60004
rect 67396 59948 67406 60004
rect 68562 59948 68572 60004
rect 68628 59948 69468 60004
rect 69524 59948 69534 60004
rect 70802 59948 70812 60004
rect 70868 59948 71932 60004
rect 71988 59948 71998 60004
rect 72594 59948 72604 60004
rect 72660 59948 74508 60004
rect 74564 59948 78092 60004
rect 78148 59948 78158 60004
rect 81666 59948 81676 60004
rect 81732 59948 82012 60004
rect 82068 59948 84364 60004
rect 84420 59948 84430 60004
rect 84802 59948 84812 60004
rect 84868 59948 85596 60004
rect 85652 59948 85662 60004
rect 86034 59948 86044 60004
rect 86100 59948 89068 60004
rect 89124 59948 89134 60004
rect 94322 59948 94332 60004
rect 94388 59948 97692 60004
rect 97748 59948 97758 60004
rect 56802 59836 56812 59892
rect 56868 59836 57260 59892
rect 57316 59836 57326 59892
rect 58034 59836 58044 59892
rect 58100 59836 58380 59892
rect 58436 59836 60508 59892
rect 60564 59836 60574 59892
rect 65090 59836 65100 59892
rect 65156 59836 66780 59892
rect 66836 59836 66846 59892
rect 76402 59836 76412 59892
rect 76468 59836 78428 59892
rect 78484 59836 78494 59892
rect 80210 59836 80220 59892
rect 80276 59836 84476 59892
rect 84532 59836 84542 59892
rect 97346 59836 97356 59892
rect 97412 59836 98028 59892
rect 98084 59836 98094 59892
rect 57362 59724 57372 59780
rect 57428 59724 58492 59780
rect 58548 59724 58558 59780
rect 65538 59724 65548 59780
rect 65604 59724 66332 59780
rect 66388 59724 68572 59780
rect 68628 59724 68638 59780
rect 70242 59724 70252 59780
rect 70308 59724 70476 59780
rect 70532 59724 77308 59780
rect 77364 59724 78204 59780
rect 78260 59724 81116 59780
rect 81172 59724 81900 59780
rect 81956 59724 81966 59780
rect 88386 59724 88396 59780
rect 88452 59724 88844 59780
rect 88900 59724 89404 59780
rect 89460 59724 89470 59780
rect 58492 59668 58548 59724
rect 54338 59612 54348 59668
rect 54404 59612 58156 59668
rect 58212 59612 58222 59668
rect 58492 59612 58940 59668
rect 58996 59612 77532 59668
rect 77588 59612 77598 59668
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 81266 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81550 59612
rect 56466 59500 56476 59556
rect 56532 59500 58492 59556
rect 58548 59500 58558 59556
rect 65426 59500 65436 59556
rect 65492 59500 68460 59556
rect 68516 59500 68526 59556
rect 70578 59500 70588 59556
rect 70644 59500 70924 59556
rect 70980 59500 73724 59556
rect 73780 59500 73790 59556
rect 82114 59500 82124 59556
rect 82180 59500 83692 59556
rect 83748 59500 83758 59556
rect 73724 59444 73780 59500
rect 47954 59388 47964 59444
rect 48020 59388 48748 59444
rect 48804 59388 49196 59444
rect 49252 59388 50428 59444
rect 50484 59388 50494 59444
rect 54450 59388 54460 59444
rect 54516 59388 58156 59444
rect 58212 59388 58222 59444
rect 61058 59388 61068 59444
rect 61124 59388 61740 59444
rect 61796 59388 63868 59444
rect 63924 59388 63934 59444
rect 73724 59388 74844 59444
rect 74900 59388 74910 59444
rect 80882 59388 80892 59444
rect 80948 59388 83468 59444
rect 83524 59388 83534 59444
rect 87490 59388 87500 59444
rect 87556 59388 89852 59444
rect 89908 59388 90244 59444
rect 47842 59276 47852 59332
rect 47908 59276 50316 59332
rect 50372 59276 50382 59332
rect 56802 59276 56812 59332
rect 56868 59276 57596 59332
rect 57652 59276 57662 59332
rect 68562 59276 68572 59332
rect 68628 59276 69356 59332
rect 69412 59276 71484 59332
rect 71540 59276 71550 59332
rect 73490 59276 73500 59332
rect 73556 59276 78988 59332
rect 79044 59276 88172 59332
rect 88228 59276 88238 59332
rect 46946 59164 46956 59220
rect 47012 59164 48524 59220
rect 48580 59164 54236 59220
rect 54292 59164 54302 59220
rect 57698 59164 57708 59220
rect 57764 59164 58940 59220
rect 58996 59164 59006 59220
rect 63970 59164 63980 59220
rect 64036 59164 65324 59220
rect 65380 59164 65390 59220
rect 79314 59164 79324 59220
rect 79380 59164 79996 59220
rect 80052 59164 80062 59220
rect 61842 59052 61852 59108
rect 61908 59052 62412 59108
rect 62468 59052 65772 59108
rect 65828 59052 65838 59108
rect 66882 59052 66892 59108
rect 66948 59052 69244 59108
rect 69300 59052 70476 59108
rect 70532 59052 70542 59108
rect 75842 59052 75852 59108
rect 75908 59052 79772 59108
rect 79828 59052 79838 59108
rect 82226 59052 82236 59108
rect 82292 59052 82572 59108
rect 82628 59052 82638 59108
rect 84466 59052 84476 59108
rect 84532 59052 85260 59108
rect 85316 59052 86380 59108
rect 86436 59052 86446 59108
rect 90188 58996 90244 59388
rect 94434 59276 94444 59332
rect 94500 59276 95564 59332
rect 95620 59276 95630 59332
rect 52434 58940 52444 58996
rect 52500 58940 57932 58996
rect 57988 58940 57998 58996
rect 62738 58940 62748 58996
rect 62804 58940 63532 58996
rect 63588 58940 63598 58996
rect 74610 58940 74620 58996
rect 74676 58940 76188 58996
rect 76244 58940 76972 58996
rect 77028 58940 82124 58996
rect 82180 58940 82190 58996
rect 90178 58940 90188 58996
rect 90244 58940 90254 58996
rect 55458 58828 55468 58884
rect 55524 58828 57260 58884
rect 57316 58828 57326 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 96626 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96910 58828
rect 71362 58716 71372 58772
rect 71428 58716 72044 58772
rect 72100 58716 72110 58772
rect 78306 58716 78316 58772
rect 78372 58716 81004 58772
rect 81060 58716 81070 58772
rect 54450 58604 54460 58660
rect 54516 58604 57596 58660
rect 57652 58604 57662 58660
rect 63186 58604 63196 58660
rect 63252 58604 64988 58660
rect 65044 58604 65054 58660
rect 69570 58604 69580 58660
rect 69636 58604 70812 58660
rect 70868 58604 70878 58660
rect 71474 58604 71484 58660
rect 71540 58604 83132 58660
rect 83188 58604 84028 58660
rect 84084 58604 84812 58660
rect 84868 58604 84878 58660
rect 50530 58492 50540 58548
rect 50596 58492 51996 58548
rect 52052 58492 67004 58548
rect 67060 58492 67070 58548
rect 68114 58492 68124 58548
rect 68180 58492 69244 58548
rect 69300 58492 70252 58548
rect 70308 58492 70318 58548
rect 74274 58492 74284 58548
rect 74340 58492 76076 58548
rect 76132 58492 78204 58548
rect 78260 58492 78270 58548
rect 78418 58492 78428 58548
rect 78484 58492 80220 58548
rect 80276 58492 80286 58548
rect 85362 58492 85372 58548
rect 85428 58492 88508 58548
rect 88564 58492 88574 58548
rect 90066 58492 90076 58548
rect 90132 58492 90636 58548
rect 90692 58492 90702 58548
rect 48514 58380 48524 58436
rect 48580 58380 49420 58436
rect 49476 58380 49486 58436
rect 55234 58380 55244 58436
rect 55300 58380 58492 58436
rect 58548 58380 59612 58436
rect 59668 58380 59836 58436
rect 59892 58380 60956 58436
rect 61012 58380 64204 58436
rect 64260 58380 64540 58436
rect 64596 58380 64606 58436
rect 65090 58380 65100 58436
rect 65156 58380 65884 58436
rect 65940 58380 65950 58436
rect 68226 58380 68236 58436
rect 68292 58380 68572 58436
rect 68628 58380 73612 58436
rect 73668 58380 74172 58436
rect 74228 58380 74238 58436
rect 75618 58380 75628 58436
rect 75684 58380 79100 58436
rect 79156 58380 79772 58436
rect 79828 58380 79838 58436
rect 91410 58380 91420 58436
rect 91476 58380 91756 58436
rect 91812 58380 91980 58436
rect 92036 58380 92046 58436
rect 54674 58268 54684 58324
rect 54740 58268 55916 58324
rect 55972 58268 55982 58324
rect 60610 58268 60620 58324
rect 60676 58268 65548 58324
rect 65604 58268 65614 58324
rect 69458 58268 69468 58324
rect 69524 58268 71596 58324
rect 71652 58268 71820 58324
rect 71876 58268 71886 58324
rect 73042 58268 73052 58324
rect 73108 58268 74060 58324
rect 74116 58268 74126 58324
rect 74610 58268 74620 58324
rect 74676 58268 77084 58324
rect 77140 58268 77150 58324
rect 77634 58268 77644 58324
rect 77700 58268 78204 58324
rect 78260 58268 81564 58324
rect 81620 58268 81630 58324
rect 84914 58268 84924 58324
rect 84980 58268 87836 58324
rect 87892 58268 89292 58324
rect 89348 58268 89358 58324
rect 94882 58268 94892 58324
rect 94948 58268 97580 58324
rect 97636 58268 97646 58324
rect 64306 58156 64316 58212
rect 64372 58156 64988 58212
rect 65044 58156 65660 58212
rect 65716 58156 65726 58212
rect 66098 58156 66108 58212
rect 66164 58156 66444 58212
rect 66500 58156 66892 58212
rect 66948 58156 66958 58212
rect 72146 58156 72156 58212
rect 72212 58156 72828 58212
rect 72884 58156 76524 58212
rect 76580 58156 77196 58212
rect 77252 58156 77262 58212
rect 78530 58156 78540 58212
rect 78596 58156 79436 58212
rect 79492 58156 79502 58212
rect 79660 58156 81676 58212
rect 81732 58156 81742 58212
rect 84476 58156 86492 58212
rect 86548 58156 87276 58212
rect 87332 58156 87342 58212
rect 72156 58100 72212 58156
rect 79660 58100 79716 58156
rect 71810 58044 71820 58100
rect 71876 58044 72212 58100
rect 74050 58044 74060 58100
rect 74116 58044 75516 58100
rect 75572 58044 77420 58100
rect 77476 58044 78876 58100
rect 78932 58044 78942 58100
rect 79314 58044 79324 58100
rect 79380 58044 79716 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 81266 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81550 58044
rect 84476 57988 84532 58156
rect 85652 58044 96460 58100
rect 96516 58044 96908 58100
rect 96964 58044 97356 58100
rect 97412 58044 97422 58100
rect 70130 57932 70140 57988
rect 70196 57932 75292 57988
rect 75348 57932 78540 57988
rect 78596 57932 80668 57988
rect 80724 57932 80734 57988
rect 84466 57932 84476 57988
rect 84532 57932 84542 57988
rect 85652 57876 85708 58044
rect 57362 57820 57372 57876
rect 57428 57820 58380 57876
rect 58436 57820 58446 57876
rect 61394 57820 61404 57876
rect 61460 57820 65548 57876
rect 65604 57820 65614 57876
rect 70354 57820 70364 57876
rect 70420 57820 73164 57876
rect 73220 57820 73230 57876
rect 74162 57820 74172 57876
rect 74228 57820 76972 57876
rect 77028 57820 78428 57876
rect 78484 57820 78494 57876
rect 78866 57820 78876 57876
rect 78932 57820 80332 57876
rect 80388 57820 82012 57876
rect 82068 57820 85708 57876
rect 92764 57820 96124 57876
rect 96180 57820 96190 57876
rect 92764 57764 92820 57820
rect 57250 57708 57260 57764
rect 57316 57708 57708 57764
rect 57764 57708 57932 57764
rect 57988 57708 57998 57764
rect 75058 57708 75068 57764
rect 75124 57708 75404 57764
rect 75460 57708 75852 57764
rect 75908 57708 76860 57764
rect 76916 57708 76926 57764
rect 77074 57708 77084 57764
rect 77140 57708 79324 57764
rect 79380 57708 79390 57764
rect 79538 57708 79548 57764
rect 79604 57708 80668 57764
rect 80724 57708 81340 57764
rect 81396 57708 81406 57764
rect 83794 57708 83804 57764
rect 83860 57708 84700 57764
rect 84756 57708 84766 57764
rect 92306 57708 92316 57764
rect 92372 57708 92764 57764
rect 92820 57708 92830 57764
rect 94322 57708 94332 57764
rect 94388 57708 95340 57764
rect 95396 57708 95406 57764
rect 77084 57652 77140 57708
rect 52994 57596 53004 57652
rect 53060 57596 57372 57652
rect 57428 57596 57438 57652
rect 72482 57596 72492 57652
rect 72548 57596 73388 57652
rect 73444 57596 73454 57652
rect 73714 57596 73724 57652
rect 73780 57596 74284 57652
rect 74340 57596 74350 57652
rect 76514 57596 76524 57652
rect 76580 57596 77140 57652
rect 85922 57596 85932 57652
rect 85988 57596 87500 57652
rect 87556 57596 87566 57652
rect 88610 57596 88620 57652
rect 88676 57596 91420 57652
rect 91476 57596 91486 57652
rect 92194 57596 92204 57652
rect 92260 57596 92428 57652
rect 92484 57596 93660 57652
rect 93716 57596 93726 57652
rect 50754 57484 50764 57540
rect 50820 57484 52220 57540
rect 52276 57484 52780 57540
rect 52836 57484 52846 57540
rect 68114 57484 68124 57540
rect 68180 57484 68796 57540
rect 68852 57484 68862 57540
rect 70578 57484 70588 57540
rect 70644 57484 70812 57540
rect 70868 57484 71372 57540
rect 71428 57484 72604 57540
rect 72660 57484 72670 57540
rect 83458 57372 83468 57428
rect 83524 57372 86828 57428
rect 86884 57372 88172 57428
rect 88228 57372 88238 57428
rect 82898 57260 82908 57316
rect 82964 57260 83916 57316
rect 83972 57260 83982 57316
rect 86930 57260 86940 57316
rect 86996 57260 87724 57316
rect 87780 57260 87948 57316
rect 88004 57260 88508 57316
rect 88564 57260 88574 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 96626 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96910 57260
rect 69682 57148 69692 57204
rect 69748 57148 70140 57204
rect 70196 57148 70206 57204
rect 74918 57148 74956 57204
rect 75012 57148 75022 57204
rect 77410 57148 77420 57204
rect 77476 57148 78316 57204
rect 78372 57148 78382 57204
rect 83794 57148 83804 57204
rect 83860 57148 87388 57204
rect 87444 57148 87454 57204
rect 88610 57148 88620 57204
rect 88676 57148 89516 57204
rect 89572 57148 89582 57204
rect 2146 57036 2156 57092
rect 2212 57036 55468 57092
rect 56690 57036 56700 57092
rect 56756 57036 57484 57092
rect 57540 57036 57550 57092
rect 60386 57036 60396 57092
rect 60452 57036 60620 57092
rect 60676 57036 64764 57092
rect 64820 57036 64830 57092
rect 71138 57036 71148 57092
rect 71204 57036 72156 57092
rect 72212 57036 72222 57092
rect 74722 57036 74732 57092
rect 74788 57036 75292 57092
rect 75348 57036 75358 57092
rect 77298 57036 77308 57092
rect 77364 57036 79996 57092
rect 80052 57036 80062 57092
rect 55412 56980 55468 57036
rect 77308 56980 77364 57036
rect 49746 56924 49756 56980
rect 49812 56924 51212 56980
rect 51268 56924 51996 56980
rect 52052 56924 52062 56980
rect 53330 56924 53340 56980
rect 53396 56924 54348 56980
rect 54404 56924 54414 56980
rect 55412 56924 70588 56980
rect 70644 56924 70654 56980
rect 74050 56924 74060 56980
rect 74116 56924 74844 56980
rect 74900 56924 77364 56980
rect 78978 56924 78988 56980
rect 79044 56924 79548 56980
rect 79604 56924 79614 56980
rect 80546 56924 80556 56980
rect 80612 56924 81116 56980
rect 81172 56924 81182 56980
rect 93090 56924 93100 56980
rect 93156 56924 95004 56980
rect 95060 56924 95070 56980
rect 57474 56812 57484 56868
rect 57540 56812 58324 56868
rect 93650 56812 93660 56868
rect 93716 56812 94332 56868
rect 94388 56812 94398 56868
rect 58268 56756 58324 56812
rect 56466 56700 56476 56756
rect 56532 56700 57372 56756
rect 57428 56700 57438 56756
rect 58258 56700 58268 56756
rect 58324 56700 58716 56756
rect 58772 56700 58782 56756
rect 66882 56700 66892 56756
rect 66948 56700 75460 56756
rect 81778 56700 81788 56756
rect 81844 56700 82348 56756
rect 82404 56700 82684 56756
rect 82740 56700 82750 56756
rect 75404 56644 75460 56700
rect 56578 56588 56588 56644
rect 56644 56588 58156 56644
rect 58212 56588 58222 56644
rect 67106 56588 67116 56644
rect 67172 56588 71148 56644
rect 71204 56588 74172 56644
rect 74228 56588 74238 56644
rect 75394 56588 75404 56644
rect 75460 56588 77420 56644
rect 77476 56588 79436 56644
rect 79492 56588 79502 56644
rect 80546 56588 80556 56644
rect 80612 56588 81452 56644
rect 81508 56588 81518 56644
rect 81890 56588 81900 56644
rect 81956 56588 82796 56644
rect 82852 56588 83020 56644
rect 83076 56588 83086 56644
rect 91858 56588 91868 56644
rect 91924 56588 93324 56644
rect 93380 56588 93390 56644
rect 93874 56588 93884 56644
rect 93940 56588 95564 56644
rect 95620 56588 95630 56644
rect 71474 56476 71484 56532
rect 71540 56476 72044 56532
rect 72100 56476 76300 56532
rect 76356 56476 77868 56532
rect 77924 56476 77934 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 81266 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81550 56476
rect 48290 56364 48300 56420
rect 48356 56364 49644 56420
rect 49700 56364 49710 56420
rect 54450 56364 54460 56420
rect 54516 56364 57596 56420
rect 57652 56364 57662 56420
rect 70914 56364 70924 56420
rect 70980 56364 72604 56420
rect 72660 56364 73948 56420
rect 74946 56364 74956 56420
rect 75012 56364 77196 56420
rect 77252 56364 77262 56420
rect 89618 56364 89628 56420
rect 89684 56364 93100 56420
rect 93156 56364 93166 56420
rect 48402 56252 48412 56308
rect 48468 56252 49532 56308
rect 49588 56252 50652 56308
rect 50708 56252 51436 56308
rect 51492 56252 52220 56308
rect 52276 56252 52668 56308
rect 52724 56252 53564 56308
rect 53620 56252 53630 56308
rect 54562 56252 54572 56308
rect 54628 56252 57372 56308
rect 57428 56252 57438 56308
rect 71922 56252 71932 56308
rect 71988 56252 72716 56308
rect 72772 56252 72940 56308
rect 72996 56252 73006 56308
rect 73892 56252 73948 56364
rect 74004 56252 77756 56308
rect 77812 56252 77822 56308
rect 80322 56252 80332 56308
rect 80388 56252 81900 56308
rect 81956 56252 81966 56308
rect 85586 56252 85596 56308
rect 85652 56252 86604 56308
rect 86660 56252 86670 56308
rect 88610 56252 88620 56308
rect 88676 56252 90076 56308
rect 90132 56252 90142 56308
rect 90514 56252 90524 56308
rect 90580 56252 92204 56308
rect 92260 56252 92270 56308
rect 63522 56140 63532 56196
rect 63588 56140 65548 56196
rect 65604 56140 65614 56196
rect 72146 56140 72156 56196
rect 72212 56140 72380 56196
rect 72436 56140 73500 56196
rect 73556 56140 73566 56196
rect 73826 56140 73836 56196
rect 73892 56140 75852 56196
rect 75908 56140 75918 56196
rect 88274 56140 88284 56196
rect 88340 56140 90300 56196
rect 90356 56140 90366 56196
rect 56466 56028 56476 56084
rect 56532 56028 58156 56084
rect 58212 56028 58222 56084
rect 59154 56028 59164 56084
rect 59220 56028 68348 56084
rect 68404 56028 68908 56084
rect 68964 56028 69356 56084
rect 69412 56028 69422 56084
rect 75730 56028 75740 56084
rect 75796 56028 76188 56084
rect 76244 56028 76254 56084
rect 76402 56028 76412 56084
rect 76468 56028 77084 56084
rect 77140 56028 77150 56084
rect 82786 56028 82796 56084
rect 82852 56028 87500 56084
rect 87556 56028 92036 56084
rect 91980 55972 92036 56028
rect 91970 55916 91980 55972
rect 92036 55916 92316 55972
rect 92372 55916 97244 55972
rect 97300 55916 97804 55972
rect 97860 55916 97870 55972
rect 66434 55804 66444 55860
rect 66500 55804 67452 55860
rect 67508 55804 67518 55860
rect 78418 55804 78428 55860
rect 78484 55804 78876 55860
rect 78932 55804 78942 55860
rect 93538 55804 93548 55860
rect 93604 55804 94332 55860
rect 94388 55804 96236 55860
rect 96292 55804 97020 55860
rect 97076 55804 97580 55860
rect 97636 55804 97646 55860
rect 68562 55692 68572 55748
rect 68628 55692 83244 55748
rect 83300 55692 83310 55748
rect 89618 55692 89628 55748
rect 89684 55692 90636 55748
rect 90692 55692 92316 55748
rect 92372 55692 93436 55748
rect 93492 55692 93502 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 96626 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96910 55692
rect 53106 55468 53116 55524
rect 53172 55468 55468 55524
rect 55524 55468 55534 55524
rect 58146 55468 58156 55524
rect 58212 55468 60620 55524
rect 60676 55468 60686 55524
rect 74946 55468 74956 55524
rect 75012 55468 75852 55524
rect 75908 55468 75918 55524
rect 50194 55356 50204 55412
rect 50260 55356 51212 55412
rect 51268 55356 51278 55412
rect 58146 55356 58156 55412
rect 58212 55356 61180 55412
rect 61236 55356 61246 55412
rect 62402 55356 62412 55412
rect 62468 55356 63980 55412
rect 64036 55356 64046 55412
rect 68114 55356 68124 55412
rect 68180 55356 73388 55412
rect 73444 55356 74844 55412
rect 74900 55356 74910 55412
rect 75730 55356 75740 55412
rect 75796 55356 76524 55412
rect 76580 55356 76590 55412
rect 82562 55356 82572 55412
rect 82628 55356 83356 55412
rect 83412 55356 83422 55412
rect 55570 55244 55580 55300
rect 55636 55244 57036 55300
rect 57092 55244 57102 55300
rect 78194 55244 78204 55300
rect 78260 55244 79772 55300
rect 79828 55244 81788 55300
rect 81844 55244 82124 55300
rect 82180 55244 83132 55300
rect 83188 55244 84028 55300
rect 84084 55244 85148 55300
rect 85204 55244 85932 55300
rect 85988 55244 85998 55300
rect 92194 55244 92204 55300
rect 92260 55244 93548 55300
rect 93604 55244 93614 55300
rect 52098 55132 52108 55188
rect 52164 55132 52444 55188
rect 52500 55132 52510 55188
rect 60834 55132 60844 55188
rect 60900 55132 61292 55188
rect 61348 55132 61358 55188
rect 61506 55132 61516 55188
rect 61572 55132 63868 55188
rect 63924 55132 64764 55188
rect 64820 55132 65660 55188
rect 65716 55132 65726 55188
rect 73892 55132 76524 55188
rect 76580 55132 77196 55188
rect 77252 55132 77262 55188
rect 85586 55132 85596 55188
rect 85652 55132 86044 55188
rect 86100 55132 86110 55188
rect 60498 55020 60508 55076
rect 60564 55020 62412 55076
rect 62468 55020 65324 55076
rect 65380 55020 65390 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 73892 54740 73948 55132
rect 83794 55020 83804 55076
rect 83860 55020 84364 55076
rect 84420 55020 84430 55076
rect 81266 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81550 54908
rect 83010 54796 83020 54852
rect 83076 54796 92316 54852
rect 92372 54796 92764 54852
rect 92820 54796 93548 54852
rect 93604 54796 93614 54852
rect 59714 54684 59724 54740
rect 59780 54684 62300 54740
rect 62356 54684 62366 54740
rect 63074 54684 63084 54740
rect 63140 54684 64316 54740
rect 64372 54684 65324 54740
rect 65380 54684 65390 54740
rect 72258 54684 72268 54740
rect 72324 54684 74060 54740
rect 74116 54684 74126 54740
rect 74946 54684 74956 54740
rect 75012 54684 77644 54740
rect 77700 54684 77710 54740
rect 87490 54684 87500 54740
rect 87556 54684 89292 54740
rect 89348 54684 89358 54740
rect 89842 54684 89852 54740
rect 89908 54684 90860 54740
rect 90916 54684 90926 54740
rect 61394 54572 61404 54628
rect 61460 54572 62076 54628
rect 62132 54572 62142 54628
rect 62850 54572 62860 54628
rect 62916 54572 64204 54628
rect 64260 54572 64270 54628
rect 69458 54572 69468 54628
rect 69524 54572 69916 54628
rect 69972 54572 70700 54628
rect 70756 54572 71148 54628
rect 71204 54572 75852 54628
rect 75908 54572 76188 54628
rect 76244 54572 76412 54628
rect 76468 54572 76478 54628
rect 76738 54572 76748 54628
rect 76804 54572 79100 54628
rect 79156 54572 79548 54628
rect 79604 54572 80948 54628
rect 82562 54572 82572 54628
rect 82628 54572 84140 54628
rect 84196 54572 84206 54628
rect 84466 54572 84476 54628
rect 84532 54572 85260 54628
rect 85316 54572 85326 54628
rect 87826 54572 87836 54628
rect 87892 54572 89516 54628
rect 89572 54572 89582 54628
rect 90290 54572 90300 54628
rect 90356 54572 90860 54628
rect 90916 54572 90926 54628
rect 91074 54572 91084 54628
rect 91140 54572 93660 54628
rect 93716 54572 93726 54628
rect 80892 54516 80948 54572
rect 50978 54460 50988 54516
rect 51044 54460 52780 54516
rect 52836 54460 52846 54516
rect 53106 54460 53116 54516
rect 53172 54460 55020 54516
rect 55076 54460 55692 54516
rect 55748 54460 61068 54516
rect 61124 54460 61852 54516
rect 61908 54460 61918 54516
rect 77746 54460 77756 54516
rect 77812 54460 80668 54516
rect 80724 54460 80734 54516
rect 80892 54460 86828 54516
rect 86884 54460 88172 54516
rect 88228 54460 90412 54516
rect 90468 54460 91196 54516
rect 91252 54460 91262 54516
rect 79202 54348 79212 54404
rect 79268 54348 80556 54404
rect 80612 54348 80622 54404
rect 83906 54348 83916 54404
rect 83972 54348 84700 54404
rect 84756 54348 84766 54404
rect 90850 54348 90860 54404
rect 90916 54348 92092 54404
rect 92148 54348 92158 54404
rect 47954 54236 47964 54292
rect 48020 54236 51772 54292
rect 51828 54236 51838 54292
rect 56018 54236 56028 54292
rect 56084 54236 56476 54292
rect 56532 54236 57372 54292
rect 57428 54236 59276 54292
rect 59332 54236 59948 54292
rect 60004 54236 60014 54292
rect 88274 54236 88284 54292
rect 88340 54236 91644 54292
rect 91700 54236 94444 54292
rect 94500 54236 95004 54292
rect 95060 54236 95564 54292
rect 95620 54236 95630 54292
rect 89506 54124 89516 54180
rect 89572 54124 90076 54180
rect 90132 54124 90142 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 96626 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96910 54124
rect 52770 54012 52780 54068
rect 52836 54012 53452 54068
rect 53508 54012 53900 54068
rect 53956 54012 55468 54068
rect 56690 54012 56700 54068
rect 56756 54012 57484 54068
rect 57540 54012 57550 54068
rect 89954 54012 89964 54068
rect 90020 54012 90300 54068
rect 90356 54012 90366 54068
rect 93622 54012 93660 54068
rect 93716 54012 93726 54068
rect 55412 53956 55468 54012
rect 55412 53900 74844 53956
rect 74900 53900 75404 53956
rect 75460 53900 75470 53956
rect 91858 53900 91868 53956
rect 91924 53900 92092 53956
rect 92148 53900 92876 53956
rect 92932 53900 93100 53956
rect 93156 53900 93166 53956
rect 60946 53788 60956 53844
rect 61012 53788 62188 53844
rect 62244 53788 62254 53844
rect 64530 53788 64540 53844
rect 64596 53788 65548 53844
rect 65604 53788 65614 53844
rect 83346 53788 83356 53844
rect 83412 53788 85708 53844
rect 89394 53788 89404 53844
rect 89460 53788 90748 53844
rect 90804 53788 91196 53844
rect 91252 53788 92204 53844
rect 92260 53788 92270 53844
rect 85652 53732 85708 53788
rect 51650 53676 51660 53732
rect 51716 53676 53004 53732
rect 53060 53676 53070 53732
rect 56354 53676 56364 53732
rect 56420 53676 57036 53732
rect 57092 53676 57484 53732
rect 57540 53676 57820 53732
rect 57876 53676 67004 53732
rect 67060 53676 67788 53732
rect 67844 53676 74396 53732
rect 74452 53676 74462 53732
rect 76402 53676 76412 53732
rect 76468 53676 78764 53732
rect 78820 53676 78830 53732
rect 85652 53676 90860 53732
rect 90916 53676 90926 53732
rect 92530 53676 92540 53732
rect 92596 53676 94780 53732
rect 94836 53676 94846 53732
rect 97682 53676 97692 53732
rect 97748 53676 98028 53732
rect 98084 53676 98094 53732
rect 94108 53620 94164 53676
rect 48178 53564 48188 53620
rect 48244 53564 49532 53620
rect 49588 53564 49598 53620
rect 64530 53564 64540 53620
rect 64596 53564 65660 53620
rect 65716 53564 66108 53620
rect 66164 53564 67228 53620
rect 71138 53564 71148 53620
rect 71204 53564 71708 53620
rect 71764 53564 73500 53620
rect 73556 53564 73566 53620
rect 76626 53564 76636 53620
rect 76692 53564 78092 53620
rect 78148 53564 78158 53620
rect 83010 53564 83020 53620
rect 83076 53564 83580 53620
rect 83636 53564 85148 53620
rect 85204 53564 85214 53620
rect 85652 53564 86380 53620
rect 86436 53564 86940 53620
rect 86996 53564 87006 53620
rect 94098 53564 94108 53620
rect 94164 53564 94174 53620
rect 50866 53452 50876 53508
rect 50932 53452 52556 53508
rect 52612 53452 52622 53508
rect 56466 53452 56476 53508
rect 56532 53452 57036 53508
rect 57092 53452 57102 53508
rect 67172 53396 67228 53564
rect 85652 53508 85708 53564
rect 68562 53452 68572 53508
rect 68628 53452 69244 53508
rect 69300 53452 69310 53508
rect 70354 53452 70364 53508
rect 70420 53452 70924 53508
rect 70980 53452 71260 53508
rect 71316 53452 72884 53508
rect 72828 53396 72884 53452
rect 73892 53452 85708 53508
rect 86034 53452 86044 53508
rect 86100 53452 87052 53508
rect 87108 53452 87118 53508
rect 73892 53396 73948 53452
rect 67172 53340 69580 53396
rect 69636 53340 70812 53396
rect 70868 53340 71820 53396
rect 71876 53340 71886 53396
rect 72828 53340 73948 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 81266 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81550 53340
rect 52098 53116 52108 53172
rect 52164 53116 52892 53172
rect 52948 53116 52958 53172
rect 60834 53116 60844 53172
rect 60900 53116 63196 53172
rect 63252 53116 63262 53172
rect 63410 53116 63420 53172
rect 63476 53116 64316 53172
rect 64372 53116 64382 53172
rect 70354 53116 70364 53172
rect 70420 53116 71148 53172
rect 71204 53116 71214 53172
rect 74722 53116 74732 53172
rect 74788 53116 75292 53172
rect 75348 53116 75358 53172
rect 77298 53116 77308 53172
rect 77364 53116 77644 53172
rect 77700 53116 77710 53172
rect 78418 53116 78428 53172
rect 78484 53116 80220 53172
rect 80276 53116 80286 53172
rect 95666 53116 95676 53172
rect 95732 53116 96908 53172
rect 96964 53116 96974 53172
rect 63522 53004 63532 53060
rect 63588 53004 64540 53060
rect 64596 53004 64606 53060
rect 67330 53004 67340 53060
rect 67396 53004 68236 53060
rect 68292 53004 68302 53060
rect 90178 53004 90188 53060
rect 90244 53004 94668 53060
rect 94724 53004 94948 53060
rect 48850 52892 48860 52948
rect 48916 52892 49532 52948
rect 49588 52892 49598 52948
rect 52994 52892 53004 52948
rect 53060 52892 55132 52948
rect 55188 52892 55198 52948
rect 60274 52892 60284 52948
rect 60340 52892 61964 52948
rect 62020 52892 62524 52948
rect 62580 52892 62590 52948
rect 72482 52892 72492 52948
rect 72548 52892 73836 52948
rect 73892 52892 75740 52948
rect 75796 52892 75806 52948
rect 76738 52892 76748 52948
rect 76804 52892 78316 52948
rect 78372 52892 79100 52948
rect 79156 52892 90076 52948
rect 90132 52892 90142 52948
rect 93986 52892 93996 52948
rect 94052 52892 94556 52948
rect 94612 52892 94622 52948
rect 94892 52836 94948 53004
rect 96114 52892 96124 52948
rect 96180 52892 97580 52948
rect 97636 52892 97646 52948
rect 72818 52780 72828 52836
rect 72884 52780 74396 52836
rect 74452 52780 74462 52836
rect 85250 52780 85260 52836
rect 85316 52780 86044 52836
rect 86100 52780 86110 52836
rect 94892 52780 97132 52836
rect 97188 52780 97198 52836
rect 94892 52724 94948 52780
rect 94882 52668 94892 52724
rect 94948 52668 94958 52724
rect 66994 52556 67004 52612
rect 67060 52556 70028 52612
rect 70084 52556 70094 52612
rect 78754 52556 78764 52612
rect 78820 52556 79100 52612
rect 79156 52556 96124 52612
rect 96180 52556 96190 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 96626 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96910 52556
rect 67106 52444 67116 52500
rect 67172 52444 68572 52500
rect 68628 52444 68638 52500
rect 82338 52444 82348 52500
rect 82404 52444 82414 52500
rect 82348 52388 82404 52444
rect 62066 52332 62076 52388
rect 62132 52332 70812 52388
rect 70868 52332 71260 52388
rect 71316 52332 73948 52388
rect 74004 52332 74014 52388
rect 82348 52332 82684 52388
rect 82740 52332 83244 52388
rect 83300 52332 83310 52388
rect 52882 52220 52892 52276
rect 52948 52220 53340 52276
rect 53396 52220 56588 52276
rect 56644 52220 56654 52276
rect 61618 52220 61628 52276
rect 61684 52220 71708 52276
rect 71764 52220 73500 52276
rect 73556 52220 73566 52276
rect 76850 52220 76860 52276
rect 76916 52220 77644 52276
rect 77700 52220 77710 52276
rect 70140 52164 70196 52220
rect 52546 52108 52556 52164
rect 52612 52108 57596 52164
rect 57652 52108 57662 52164
rect 62626 52108 62636 52164
rect 62692 52108 63980 52164
rect 64036 52108 68572 52164
rect 68628 52108 69132 52164
rect 69188 52108 69198 52164
rect 70130 52108 70140 52164
rect 70196 52108 70206 52164
rect 85474 52108 85484 52164
rect 85540 52108 87500 52164
rect 87556 52108 87566 52164
rect 94322 52108 94332 52164
rect 94388 52108 95340 52164
rect 95396 52108 95406 52164
rect 54348 51940 54404 52108
rect 67788 52052 67844 52108
rect 67778 51996 67788 52052
rect 67844 51996 67854 52052
rect 70690 51996 70700 52052
rect 70756 51996 74060 52052
rect 74116 51996 74126 52052
rect 74722 51996 74732 52052
rect 74788 51996 74956 52052
rect 75012 51996 75022 52052
rect 90692 51996 91756 52052
rect 91812 51996 91822 52052
rect 70700 51940 70756 51996
rect 90692 51940 90748 51996
rect 54338 51884 54348 51940
rect 54404 51884 54414 51940
rect 55010 51884 55020 51940
rect 55076 51884 58268 51940
rect 58324 51884 58940 51940
rect 58996 51884 60844 51940
rect 60900 51884 60910 51940
rect 63746 51884 63756 51940
rect 63812 51884 70756 51940
rect 73714 51884 73724 51940
rect 73780 51884 75516 51940
rect 75572 51884 77420 51940
rect 77476 51884 77486 51940
rect 85698 51884 85708 51940
rect 85764 51884 86380 51940
rect 86436 51884 86446 51940
rect 86930 51884 86940 51940
rect 86996 51884 89628 51940
rect 89684 51884 90748 51940
rect 96226 51884 96236 51940
rect 96292 51884 97804 51940
rect 97860 51884 97870 51940
rect 90178 51772 90188 51828
rect 90244 51772 93660 51828
rect 93716 51772 94108 51828
rect 94164 51772 94174 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 81266 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81550 51772
rect 54114 51660 54124 51716
rect 54180 51660 55356 51716
rect 55412 51660 55422 51716
rect 58706 51548 58716 51604
rect 58772 51548 58782 51604
rect 64082 51548 64092 51604
rect 64148 51548 64764 51604
rect 64820 51548 65324 51604
rect 65380 51548 65390 51604
rect 74498 51548 74508 51604
rect 74564 51548 75068 51604
rect 75124 51548 93212 51604
rect 93268 51548 93996 51604
rect 94052 51548 94062 51604
rect 94658 51548 94668 51604
rect 94724 51548 97468 51604
rect 97524 51548 97534 51604
rect 58716 51492 58772 51548
rect 56242 51436 56252 51492
rect 56308 51436 56924 51492
rect 56980 51436 59388 51492
rect 59444 51436 59724 51492
rect 59780 51436 62076 51492
rect 62132 51436 62142 51492
rect 72034 51436 72044 51492
rect 72100 51436 73500 51492
rect 73556 51436 73948 51492
rect 74004 51436 74014 51492
rect 74508 51380 74564 51548
rect 78306 51436 78316 51492
rect 78372 51436 79436 51492
rect 79492 51436 79502 51492
rect 79986 51436 79996 51492
rect 80052 51436 81228 51492
rect 81284 51436 81294 51492
rect 81442 51436 81452 51492
rect 81508 51436 81900 51492
rect 81956 51436 82236 51492
rect 82292 51436 82302 51492
rect 94994 51436 95004 51492
rect 95060 51436 96236 51492
rect 96292 51436 97692 51492
rect 97748 51436 97758 51492
rect 79436 51380 79492 51436
rect 58706 51324 58716 51380
rect 58772 51324 60284 51380
rect 60340 51324 60350 51380
rect 60834 51324 60844 51380
rect 60900 51324 61628 51380
rect 61684 51324 61694 51380
rect 64082 51324 64092 51380
rect 64148 51324 64540 51380
rect 64596 51324 64606 51380
rect 72258 51324 72268 51380
rect 72324 51324 73276 51380
rect 73332 51324 73342 51380
rect 73602 51324 73612 51380
rect 73668 51324 74564 51380
rect 77074 51324 77084 51380
rect 77140 51324 78204 51380
rect 78260 51324 78270 51380
rect 79436 51324 79884 51380
rect 79940 51324 79950 51380
rect 61170 51212 61180 51268
rect 61236 51212 62972 51268
rect 63028 51212 63038 51268
rect 84914 51212 84924 51268
rect 84980 51212 89964 51268
rect 90020 51212 90030 51268
rect 57362 51100 57372 51156
rect 57428 51100 61740 51156
rect 61796 51100 61806 51156
rect 73602 51100 73612 51156
rect 73668 51100 75068 51156
rect 75124 51100 75134 51156
rect 81554 51100 81564 51156
rect 81620 51100 82012 51156
rect 82068 51100 93996 51156
rect 94052 51100 94062 51156
rect 59154 50988 59164 51044
rect 59220 50988 62412 51044
rect 62468 50988 62478 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 96626 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96910 50988
rect 56354 50764 56364 50820
rect 56420 50764 58828 50820
rect 58884 50764 59724 50820
rect 59780 50764 59790 50820
rect 52322 50652 52332 50708
rect 52388 50652 52398 50708
rect 53666 50652 53676 50708
rect 53732 50652 54908 50708
rect 54964 50652 54974 50708
rect 56802 50652 56812 50708
rect 56868 50652 58380 50708
rect 58436 50652 60172 50708
rect 60228 50652 60238 50708
rect 90066 50652 90076 50708
rect 90132 50652 91868 50708
rect 91924 50652 91934 50708
rect 52332 50596 52388 50652
rect 50978 50540 50988 50596
rect 51044 50540 51548 50596
rect 51604 50540 52388 50596
rect 54338 50540 54348 50596
rect 54404 50540 57484 50596
rect 57540 50540 57550 50596
rect 58034 50540 58044 50596
rect 58100 50540 58940 50596
rect 58996 50540 59006 50596
rect 67330 50540 67340 50596
rect 67396 50540 68572 50596
rect 68628 50540 70700 50596
rect 70756 50540 71148 50596
rect 71204 50540 73612 50596
rect 73668 50540 73678 50596
rect 74610 50540 74620 50596
rect 74676 50540 75852 50596
rect 75908 50540 75918 50596
rect 79538 50540 79548 50596
rect 79604 50540 82796 50596
rect 82852 50540 83804 50596
rect 83860 50540 83870 50596
rect 84802 50540 84812 50596
rect 84868 50540 91084 50596
rect 91140 50540 92428 50596
rect 92484 50540 92988 50596
rect 93044 50540 93054 50596
rect 50418 50428 50428 50484
rect 50484 50428 52332 50484
rect 52388 50428 52398 50484
rect 57586 50428 57596 50484
rect 57652 50428 58716 50484
rect 58772 50428 58782 50484
rect 62626 50428 62636 50484
rect 62692 50428 63196 50484
rect 63252 50428 63262 50484
rect 64530 50428 64540 50484
rect 64596 50428 65324 50484
rect 65380 50428 66444 50484
rect 66500 50428 66510 50484
rect 73714 50428 73724 50484
rect 73780 50428 74956 50484
rect 75012 50428 76860 50484
rect 76916 50428 77196 50484
rect 77252 50428 77262 50484
rect 81666 50428 81676 50484
rect 81732 50428 85260 50484
rect 85316 50428 85326 50484
rect 89058 50428 89068 50484
rect 89124 50428 89292 50484
rect 89348 50428 89358 50484
rect 90178 50428 90188 50484
rect 90244 50428 91532 50484
rect 91588 50428 91598 50484
rect 91858 50428 91868 50484
rect 91924 50428 92540 50484
rect 92596 50428 93884 50484
rect 93940 50428 93950 50484
rect 89292 50372 89348 50428
rect 51874 50316 51884 50372
rect 51940 50316 53004 50372
rect 53060 50316 53564 50372
rect 53620 50316 53630 50372
rect 54562 50316 54572 50372
rect 54628 50316 55076 50372
rect 65426 50316 65436 50372
rect 65492 50316 65996 50372
rect 66052 50316 66062 50372
rect 70466 50316 70476 50372
rect 70532 50316 71708 50372
rect 71764 50316 74284 50372
rect 74340 50316 74350 50372
rect 75170 50316 75180 50372
rect 75236 50316 76748 50372
rect 76804 50316 77084 50372
rect 77140 50316 77150 50372
rect 77634 50316 77644 50372
rect 77700 50316 81564 50372
rect 81620 50316 81630 50372
rect 85810 50316 85820 50372
rect 85876 50316 87276 50372
rect 87332 50316 87342 50372
rect 89292 50316 90076 50372
rect 90132 50316 90142 50372
rect 91186 50316 91196 50372
rect 91252 50316 93324 50372
rect 93380 50316 93390 50372
rect 94322 50316 94332 50372
rect 94388 50316 96348 50372
rect 96404 50316 96414 50372
rect 55020 50260 55076 50316
rect 55010 50204 55020 50260
rect 55076 50204 55086 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 74284 50148 74340 50316
rect 76178 50204 76188 50260
rect 76244 50204 79100 50260
rect 79156 50204 79166 50260
rect 94098 50204 94108 50260
rect 94164 50204 94892 50260
rect 94948 50204 94958 50260
rect 81266 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81550 50204
rect 72482 50092 72492 50148
rect 72548 50092 73388 50148
rect 73444 50092 73454 50148
rect 74284 50092 75180 50148
rect 75236 50092 75246 50148
rect 75954 50092 75964 50148
rect 76020 50092 78764 50148
rect 78820 50092 80556 50148
rect 80612 50092 80622 50148
rect 82338 50092 82348 50148
rect 82404 50092 84588 50148
rect 84644 50092 84654 50148
rect 95442 50092 95452 50148
rect 95508 50092 97468 50148
rect 97524 50092 97534 50148
rect 48066 49980 48076 50036
rect 48132 49980 56476 50036
rect 56532 49980 56542 50036
rect 56690 49980 56700 50036
rect 56756 49980 57036 50036
rect 57092 49980 57102 50036
rect 70018 49980 70028 50036
rect 70084 49980 72156 50036
rect 72212 49980 72222 50036
rect 75618 49980 75628 50036
rect 75684 49980 76412 50036
rect 76468 49980 84812 50036
rect 84868 49980 84878 50036
rect 88274 49980 88284 50036
rect 88340 49980 91196 50036
rect 91252 49980 91262 50036
rect 95666 49980 95676 50036
rect 95732 49980 96124 50036
rect 96180 49980 96190 50036
rect 52658 49868 52668 49924
rect 52724 49868 54404 49924
rect 55122 49868 55132 49924
rect 55188 49868 55580 49924
rect 55636 49868 56028 49924
rect 56084 49868 61964 49924
rect 62020 49868 62030 49924
rect 66322 49868 66332 49924
rect 66388 49868 66892 49924
rect 66948 49868 66958 49924
rect 68226 49868 68236 49924
rect 68292 49868 68908 49924
rect 68964 49868 73388 49924
rect 73444 49868 73454 49924
rect 75506 49868 75516 49924
rect 75572 49868 78428 49924
rect 78484 49868 78494 49924
rect 86482 49868 86492 49924
rect 86548 49868 90300 49924
rect 90356 49868 90748 49924
rect 90804 49868 90814 49924
rect 94882 49868 94892 49924
rect 94948 49868 95452 49924
rect 95508 49868 95518 49924
rect 95778 49868 95788 49924
rect 95844 49868 97356 49924
rect 97412 49868 97422 49924
rect 54348 49812 54404 49868
rect 95452 49812 95508 49868
rect 54338 49756 54348 49812
rect 54404 49756 54414 49812
rect 55412 49756 57484 49812
rect 57540 49756 58604 49812
rect 58660 49756 58670 49812
rect 62514 49756 62524 49812
rect 62580 49756 65324 49812
rect 65380 49756 65390 49812
rect 68002 49756 68012 49812
rect 68068 49756 68684 49812
rect 68740 49756 68750 49812
rect 69682 49756 69692 49812
rect 69748 49756 70364 49812
rect 70420 49756 70430 49812
rect 82226 49756 82236 49812
rect 82292 49756 83804 49812
rect 83860 49756 83870 49812
rect 84354 49756 84364 49812
rect 84420 49756 85036 49812
rect 85092 49756 85102 49812
rect 87266 49756 87276 49812
rect 87332 49756 87500 49812
rect 87556 49756 87566 49812
rect 87826 49756 87836 49812
rect 87892 49756 88284 49812
rect 88340 49756 88350 49812
rect 88946 49756 88956 49812
rect 89012 49756 89292 49812
rect 89348 49756 92652 49812
rect 92708 49756 92718 49812
rect 95452 49756 95676 49812
rect 95732 49756 97916 49812
rect 97972 49756 97982 49812
rect 55412 49588 55468 49756
rect 64642 49644 64652 49700
rect 64708 49644 65436 49700
rect 65492 49644 65502 49700
rect 79202 49644 79212 49700
rect 79268 49644 80444 49700
rect 80500 49644 80510 49700
rect 83570 49644 83580 49700
rect 83636 49644 85260 49700
rect 85316 49644 85326 49700
rect 85586 49644 85596 49700
rect 85652 49644 86996 49700
rect 91746 49644 91756 49700
rect 91812 49644 94780 49700
rect 94836 49644 95340 49700
rect 95396 49644 95406 49700
rect 85596 49588 85652 49644
rect 86940 49588 86996 49644
rect 54450 49532 54460 49588
rect 54516 49532 55468 49588
rect 56466 49532 56476 49588
rect 56532 49532 57484 49588
rect 57540 49532 58156 49588
rect 58212 49532 58222 49588
rect 66434 49532 66444 49588
rect 66500 49532 67452 49588
rect 67508 49532 75068 49588
rect 75124 49532 75134 49588
rect 80546 49532 80556 49588
rect 80612 49532 83020 49588
rect 83076 49532 84140 49588
rect 84196 49532 85652 49588
rect 86930 49532 86940 49588
rect 86996 49532 87006 49588
rect 87826 49532 87836 49588
rect 87892 49532 88396 49588
rect 88452 49532 88462 49588
rect 49858 49420 49868 49476
rect 49924 49420 51884 49476
rect 51940 49420 52556 49476
rect 52612 49420 52622 49476
rect 70578 49420 70588 49476
rect 70644 49420 70812 49476
rect 70868 49420 83916 49476
rect 83972 49420 84364 49476
rect 84420 49420 85820 49476
rect 85876 49420 85886 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 96626 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96910 49420
rect 68460 49308 71484 49364
rect 71540 49308 71932 49364
rect 71988 49308 71998 49364
rect 68460 49252 68516 49308
rect 58594 49196 58604 49252
rect 58660 49196 68516 49252
rect 68674 49196 68684 49252
rect 68740 49196 69916 49252
rect 69972 49196 69982 49252
rect 52658 49084 52668 49140
rect 52724 49084 54124 49140
rect 54180 49084 54190 49140
rect 75170 49084 75180 49140
rect 75236 49084 76188 49140
rect 76244 49084 76254 49140
rect 77970 49084 77980 49140
rect 78036 49084 78428 49140
rect 78484 49084 89068 49140
rect 89124 49084 89134 49140
rect 67218 48972 67228 49028
rect 67284 48972 68796 49028
rect 68852 48972 69580 49028
rect 69636 48972 69646 49028
rect 77298 48972 77308 49028
rect 77364 48972 77756 49028
rect 77812 48972 77822 49028
rect 78642 48972 78652 49028
rect 78708 48972 79100 49028
rect 79156 48972 81676 49028
rect 81732 48972 81742 49028
rect 84354 48972 84364 49028
rect 84420 48972 85596 49028
rect 85652 48972 85662 49028
rect 85922 48972 85932 49028
rect 85988 48972 86380 49028
rect 86436 48972 86446 49028
rect 61842 48860 61852 48916
rect 61908 48860 65212 48916
rect 65268 48860 65278 48916
rect 67442 48860 67452 48916
rect 67508 48860 68236 48916
rect 68292 48860 68302 48916
rect 83794 48860 83804 48916
rect 83860 48860 84588 48916
rect 84644 48860 84654 48916
rect 85026 48860 85036 48916
rect 85092 48860 85708 48916
rect 85764 48860 86268 48916
rect 86324 48860 86334 48916
rect 93762 48860 93772 48916
rect 93828 48860 95228 48916
rect 95284 48860 95294 48916
rect 50418 48748 50428 48804
rect 50484 48748 53340 48804
rect 53396 48748 53406 48804
rect 53554 48748 53564 48804
rect 53620 48748 54908 48804
rect 54964 48748 54974 48804
rect 57026 48748 57036 48804
rect 57092 48748 57596 48804
rect 57652 48748 60620 48804
rect 60676 48748 62188 48804
rect 62244 48748 62636 48804
rect 62692 48748 62702 48804
rect 75394 48748 75404 48804
rect 75460 48748 75470 48804
rect 83010 48748 83020 48804
rect 83076 48748 89292 48804
rect 89348 48748 89358 48804
rect 75404 48692 75460 48748
rect 62738 48636 62748 48692
rect 62804 48636 66892 48692
rect 66948 48636 66958 48692
rect 71250 48636 71260 48692
rect 71316 48636 75460 48692
rect 76514 48636 76524 48692
rect 76580 48636 77644 48692
rect 77700 48636 77710 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 81266 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81550 48636
rect 52770 48524 52780 48580
rect 52836 48524 54796 48580
rect 54852 48524 54862 48580
rect 62514 48524 62524 48580
rect 62580 48524 64932 48580
rect 65090 48524 65100 48580
rect 65156 48524 66332 48580
rect 66388 48524 66398 48580
rect 74946 48524 74956 48580
rect 75012 48524 75404 48580
rect 75460 48524 75470 48580
rect 64876 48468 64932 48524
rect 52434 48412 52444 48468
rect 52500 48412 53452 48468
rect 53508 48412 53900 48468
rect 53956 48412 53966 48468
rect 56578 48412 56588 48468
rect 56644 48412 58604 48468
rect 58660 48412 58670 48468
rect 61730 48412 61740 48468
rect 61796 48412 64204 48468
rect 64260 48412 64270 48468
rect 64876 48412 66948 48468
rect 67106 48412 67116 48468
rect 67172 48412 67340 48468
rect 67396 48412 72380 48468
rect 72436 48412 72716 48468
rect 72772 48412 74284 48468
rect 74340 48412 74350 48468
rect 76514 48412 76524 48468
rect 76580 48412 78092 48468
rect 78148 48412 78158 48468
rect 78306 48412 78316 48468
rect 78372 48412 80108 48468
rect 80164 48412 80174 48468
rect 52210 48300 52220 48356
rect 52276 48300 54124 48356
rect 54180 48300 54190 48356
rect 56466 48300 56476 48356
rect 56532 48300 57372 48356
rect 57428 48300 57438 48356
rect 62850 48300 62860 48356
rect 62916 48300 65548 48356
rect 65604 48300 65614 48356
rect 53666 48188 53676 48244
rect 53732 48188 54908 48244
rect 54964 48188 54974 48244
rect 56578 48188 56588 48244
rect 56644 48188 58380 48244
rect 58436 48188 58940 48244
rect 58996 48188 59006 48244
rect 60610 48188 60620 48244
rect 60676 48188 63476 48244
rect 64306 48188 64316 48244
rect 64372 48188 65884 48244
rect 65940 48188 66108 48244
rect 66164 48188 66174 48244
rect 63420 48132 63476 48188
rect 66892 48132 66948 48412
rect 71586 48300 71596 48356
rect 71652 48300 72268 48356
rect 72324 48300 72334 48356
rect 82338 48300 82348 48356
rect 82404 48300 82796 48356
rect 82852 48300 82862 48356
rect 92194 48300 92204 48356
rect 92260 48300 92876 48356
rect 92932 48300 92942 48356
rect 96226 48300 96236 48356
rect 96292 48300 97468 48356
rect 97524 48300 97534 48356
rect 76738 48188 76748 48244
rect 76804 48188 77532 48244
rect 77588 48188 78652 48244
rect 78708 48188 78718 48244
rect 93650 48188 93660 48244
rect 93716 48188 94220 48244
rect 94276 48188 94780 48244
rect 94836 48188 94846 48244
rect 97244 48132 97300 48300
rect 52658 48076 52668 48132
rect 52724 48076 53564 48132
rect 53620 48076 53630 48132
rect 55234 48076 55244 48132
rect 55300 48076 55692 48132
rect 55748 48076 57708 48132
rect 57764 48076 59724 48132
rect 59780 48076 62188 48132
rect 63410 48076 63420 48132
rect 63476 48076 65436 48132
rect 65492 48076 65502 48132
rect 66882 48076 66892 48132
rect 66948 48076 67452 48132
rect 67508 48076 67518 48132
rect 73826 48076 73836 48132
rect 73892 48076 78092 48132
rect 78148 48076 78158 48132
rect 86482 48076 86492 48132
rect 86548 48076 88620 48132
rect 88676 48076 90748 48132
rect 93426 48076 93436 48132
rect 93492 48076 94332 48132
rect 94388 48076 94398 48132
rect 97234 48076 97244 48132
rect 97300 48076 97310 48132
rect 60834 47964 60844 48020
rect 60900 47964 61852 48020
rect 61908 47964 61918 48020
rect 62132 47908 62188 48076
rect 90692 48020 90748 48076
rect 62290 47964 62300 48020
rect 62356 47964 64204 48020
rect 64260 47964 64270 48020
rect 65772 47964 67900 48020
rect 67956 47964 69356 48020
rect 69412 47964 69422 48020
rect 87714 47964 87724 48020
rect 87780 47964 88060 48020
rect 88116 47964 88126 48020
rect 90692 47964 94444 48020
rect 94500 47964 94510 48020
rect 94668 47964 98252 48020
rect 98308 47964 98318 48020
rect 65772 47908 65828 47964
rect 94668 47908 94724 47964
rect 62132 47852 65828 47908
rect 66882 47852 66892 47908
rect 66948 47852 68684 47908
rect 68740 47852 68750 47908
rect 90692 47852 94724 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 55234 47740 55244 47796
rect 55300 47740 59276 47796
rect 59332 47740 59342 47796
rect 73042 47628 73052 47684
rect 73108 47628 73612 47684
rect 73668 47628 73678 47684
rect 81004 47628 81788 47684
rect 81844 47628 85148 47684
rect 85204 47628 85820 47684
rect 85876 47628 88172 47684
rect 88228 47628 88238 47684
rect 81004 47572 81060 47628
rect 50082 47516 50092 47572
rect 50148 47516 53116 47572
rect 53172 47516 53182 47572
rect 55412 47516 59948 47572
rect 60004 47516 61404 47572
rect 61460 47516 61852 47572
rect 61908 47516 61918 47572
rect 77634 47516 77644 47572
rect 77700 47516 81004 47572
rect 81060 47516 81070 47572
rect 81666 47516 81676 47572
rect 81732 47516 82236 47572
rect 82292 47516 84476 47572
rect 84532 47516 84542 47572
rect 55412 47460 55468 47516
rect 54898 47404 54908 47460
rect 54964 47404 55468 47460
rect 60610 47404 60620 47460
rect 60676 47404 61516 47460
rect 61572 47404 61582 47460
rect 66098 47404 66108 47460
rect 66164 47404 66556 47460
rect 66612 47404 67004 47460
rect 67060 47404 67070 47460
rect 69570 47404 69580 47460
rect 69636 47404 70812 47460
rect 70868 47404 70878 47460
rect 76402 47404 76412 47460
rect 76468 47404 77196 47460
rect 77252 47404 77262 47460
rect 85474 47404 85484 47460
rect 85540 47404 87724 47460
rect 87780 47404 87790 47460
rect 90692 47348 90748 47852
rect 96626 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96910 47852
rect 94882 47740 94892 47796
rect 94948 47740 96236 47796
rect 96292 47740 96302 47796
rect 90962 47516 90972 47572
rect 91028 47516 92092 47572
rect 92148 47516 92158 47572
rect 93538 47404 93548 47460
rect 93604 47404 94220 47460
rect 94276 47404 95564 47460
rect 95620 47404 95630 47460
rect 96450 47404 96460 47460
rect 96516 47404 97580 47460
rect 97636 47404 97646 47460
rect 61058 47292 61068 47348
rect 61124 47292 61404 47348
rect 61460 47292 61964 47348
rect 62020 47292 62524 47348
rect 62580 47292 62590 47348
rect 64652 47292 68180 47348
rect 68338 47292 68348 47348
rect 68404 47292 68572 47348
rect 68628 47292 70028 47348
rect 70084 47292 70094 47348
rect 72258 47292 72268 47348
rect 72324 47292 72828 47348
rect 72884 47292 73388 47348
rect 73444 47292 74732 47348
rect 74788 47292 90748 47348
rect 93202 47292 93212 47348
rect 93268 47292 93660 47348
rect 93716 47292 94108 47348
rect 94164 47292 95228 47348
rect 95284 47292 95294 47348
rect 64652 47236 64708 47292
rect 68124 47236 68180 47292
rect 62132 47180 64708 47236
rect 64866 47180 64876 47236
rect 64932 47180 65660 47236
rect 65716 47180 66220 47236
rect 66276 47180 66286 47236
rect 68124 47180 70364 47236
rect 70420 47180 71260 47236
rect 71316 47180 71326 47236
rect 86034 47180 86044 47236
rect 86100 47180 87612 47236
rect 87668 47180 87678 47236
rect 88498 47180 88508 47236
rect 88564 47180 89740 47236
rect 89796 47180 89806 47236
rect 93314 47180 93324 47236
rect 93380 47180 94556 47236
rect 94612 47180 94622 47236
rect 62132 47124 62188 47180
rect 53330 47068 53340 47124
rect 53396 47068 53676 47124
rect 53732 47068 53742 47124
rect 58258 47068 58268 47124
rect 58324 47068 59052 47124
rect 59108 47068 59118 47124
rect 59490 47068 59500 47124
rect 59556 47068 62188 47124
rect 64194 47068 64204 47124
rect 64260 47068 66332 47124
rect 66388 47068 66398 47124
rect 68450 47068 68460 47124
rect 68516 47068 69244 47124
rect 69300 47068 69310 47124
rect 89842 47068 89852 47124
rect 89908 47068 93996 47124
rect 94052 47068 94062 47124
rect 94210 47068 94220 47124
rect 94276 47068 94314 47124
rect 94444 47068 96796 47124
rect 96852 47068 96862 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 81266 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81550 47068
rect 94444 47012 94500 47068
rect 93874 46956 93884 47012
rect 93940 46956 94332 47012
rect 94388 46956 94500 47012
rect 53666 46844 53676 46900
rect 53732 46844 54236 46900
rect 54292 46844 55244 46900
rect 55300 46844 55310 46900
rect 70578 46844 70588 46900
rect 70644 46844 73164 46900
rect 73220 46844 73230 46900
rect 73938 46844 73948 46900
rect 74004 46844 75852 46900
rect 75908 46844 76300 46900
rect 76356 46844 76366 46900
rect 82562 46844 82572 46900
rect 82628 46844 83132 46900
rect 83188 46844 83198 46900
rect 91410 46844 91420 46900
rect 91476 46844 91980 46900
rect 92036 46844 93772 46900
rect 93828 46844 93838 46900
rect 95554 46844 95564 46900
rect 95620 46844 96012 46900
rect 96068 46844 96078 46900
rect 60946 46732 60956 46788
rect 61012 46732 62188 46788
rect 62244 46732 62254 46788
rect 64306 46732 64316 46788
rect 64372 46732 65548 46788
rect 65604 46732 65614 46788
rect 72482 46732 72492 46788
rect 72548 46732 73836 46788
rect 73892 46732 73902 46788
rect 75058 46732 75068 46788
rect 75124 46732 75516 46788
rect 75572 46732 75582 46788
rect 85586 46732 85596 46788
rect 85652 46732 86268 46788
rect 86324 46732 86334 46788
rect 69682 46508 69692 46564
rect 69748 46508 70140 46564
rect 70196 46508 70206 46564
rect 80994 46508 81004 46564
rect 81060 46508 81676 46564
rect 81732 46508 82236 46564
rect 82292 46508 93660 46564
rect 93716 46508 93726 46564
rect 93090 46396 93100 46452
rect 93156 46396 95116 46452
rect 95172 46396 97356 46452
rect 97412 46396 97422 46452
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 73154 45948 73164 46004
rect 73220 45948 76076 46004
rect 76132 45948 76142 46004
rect 88610 45948 88620 46004
rect 88676 45948 89068 46004
rect 89124 45948 90748 46004
rect 90850 45948 90860 46004
rect 90916 45948 91308 46004
rect 91364 45948 92428 46004
rect 92484 45948 92988 46004
rect 93044 45948 93054 46004
rect 90692 45892 90748 45948
rect 82562 45836 82572 45892
rect 82628 45836 84252 45892
rect 84308 45836 85708 45892
rect 85764 45836 85774 45892
rect 89730 45836 89740 45892
rect 89796 45836 90524 45892
rect 90580 45836 90590 45892
rect 90692 45836 91196 45892
rect 91252 45836 93324 45892
rect 93380 45836 93390 45892
rect 77410 45724 77420 45780
rect 77476 45724 79100 45780
rect 79156 45724 79166 45780
rect 80658 45724 80668 45780
rect 80724 45724 82796 45780
rect 82852 45724 84476 45780
rect 84532 45724 85932 45780
rect 85988 45724 85998 45780
rect 86258 45724 86268 45780
rect 86324 45724 87724 45780
rect 87780 45724 87790 45780
rect 90738 45724 90748 45780
rect 90804 45724 92540 45780
rect 92596 45724 92606 45780
rect 80668 45668 80724 45724
rect 77858 45612 77868 45668
rect 77924 45612 79212 45668
rect 79268 45612 80724 45668
rect 83346 45612 83356 45668
rect 83412 45612 84924 45668
rect 84980 45612 84990 45668
rect 89618 45612 89628 45668
rect 89684 45612 91980 45668
rect 92036 45612 93100 45668
rect 93156 45612 93166 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 63522 45388 63532 45444
rect 63588 45388 65324 45444
rect 65380 45388 65390 45444
rect 52882 45276 52892 45332
rect 52948 45276 54124 45332
rect 54180 45276 55468 45332
rect 55524 45276 56700 45332
rect 56756 45276 56766 45332
rect 66994 45052 67004 45108
rect 67060 45052 67452 45108
rect 67508 45052 69468 45108
rect 69524 45052 70140 45108
rect 70196 45052 72268 45108
rect 72324 45052 72334 45108
rect 77186 45052 77196 45108
rect 77252 45052 77756 45108
rect 77812 45052 80668 45108
rect 80724 45052 81116 45108
rect 81172 45052 81340 45108
rect 81396 45052 81406 45108
rect 61394 44940 61404 44996
rect 61460 44940 66444 44996
rect 66500 44940 66510 44996
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 75058 44604 75068 44660
rect 75124 44604 76076 44660
rect 76132 44604 76142 44660
rect 58146 44492 58156 44548
rect 58212 44492 58492 44548
rect 58548 44492 58828 44548
rect 58884 44492 59276 44548
rect 59332 44492 59342 44548
rect 56690 44380 56700 44436
rect 56756 44380 58604 44436
rect 58660 44380 58670 44436
rect 71250 44380 71260 44436
rect 71316 44380 72380 44436
rect 72436 44380 72446 44436
rect 74386 44380 74396 44436
rect 74452 44380 75628 44436
rect 75684 44380 75694 44436
rect 75954 44380 75964 44436
rect 76020 44380 76524 44436
rect 76580 44380 77756 44436
rect 77812 44380 77822 44436
rect 95778 44380 95788 44436
rect 95844 44380 95854 44436
rect 91970 44268 91980 44324
rect 92036 44268 93548 44324
rect 93604 44268 93614 44324
rect 48738 44156 48748 44212
rect 48804 44156 49756 44212
rect 49812 44156 49822 44212
rect 61842 44156 61852 44212
rect 61908 44156 67228 44212
rect 67284 44156 67294 44212
rect 78530 44156 78540 44212
rect 78596 44156 80444 44212
rect 80500 44156 80510 44212
rect 49074 44044 49084 44100
rect 49140 44044 50092 44100
rect 50148 44044 52332 44100
rect 52388 44044 53228 44100
rect 53284 44044 53294 44100
rect 72258 44044 72268 44100
rect 72324 44044 72828 44100
rect 72884 44044 72894 44100
rect 90066 44044 90076 44100
rect 90132 44044 90636 44100
rect 90692 44044 91308 44100
rect 91364 44044 91374 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 95788 43876 95844 44380
rect 59602 43820 59612 43876
rect 59668 43820 68012 43876
rect 68068 43820 68078 43876
rect 95788 43820 95900 43876
rect 95956 43820 95966 43876
rect 62514 43708 62524 43764
rect 62580 43708 63420 43764
rect 63476 43708 63486 43764
rect 72370 43708 72380 43764
rect 72436 43708 77756 43764
rect 77812 43708 77822 43764
rect 95778 43708 95788 43764
rect 95844 43708 96236 43764
rect 96292 43708 97020 43764
rect 97076 43708 97086 43764
rect 52770 43596 52780 43652
rect 52836 43596 54348 43652
rect 54404 43596 54414 43652
rect 56578 43596 56588 43652
rect 56644 43596 57596 43652
rect 57652 43596 57662 43652
rect 64194 43596 64204 43652
rect 64260 43596 66332 43652
rect 66388 43596 66398 43652
rect 72034 43596 72044 43652
rect 72100 43596 72716 43652
rect 72772 43596 72782 43652
rect 77074 43596 77084 43652
rect 77140 43596 77868 43652
rect 77924 43596 77934 43652
rect 95554 43596 95564 43652
rect 95620 43596 97692 43652
rect 97748 43596 97758 43652
rect 48514 43484 48524 43540
rect 48580 43484 49756 43540
rect 49812 43484 49822 43540
rect 50866 43484 50876 43540
rect 50932 43484 52220 43540
rect 52276 43484 53452 43540
rect 53508 43484 53788 43540
rect 53844 43484 55468 43540
rect 64530 43484 64540 43540
rect 64596 43484 65324 43540
rect 65380 43484 65390 43540
rect 65762 43484 65772 43540
rect 65828 43484 66780 43540
rect 66836 43484 66846 43540
rect 70018 43484 70028 43540
rect 70084 43484 70924 43540
rect 70980 43484 70990 43540
rect 91410 43484 91420 43540
rect 91476 43484 92652 43540
rect 92708 43484 92718 43540
rect 55412 43428 55468 43484
rect 50082 43372 50092 43428
rect 50148 43372 51996 43428
rect 52052 43372 52062 43428
rect 55412 43372 58716 43428
rect 58772 43372 59276 43428
rect 59332 43372 69356 43428
rect 69412 43372 70364 43428
rect 70420 43372 71484 43428
rect 71540 43372 71550 43428
rect 50754 43260 50764 43316
rect 50820 43260 52332 43316
rect 52388 43260 53340 43316
rect 53396 43260 53406 43316
rect 60386 43260 60396 43316
rect 60452 43260 62076 43316
rect 62132 43260 62142 43316
rect 64418 43260 64428 43316
rect 64484 43260 65772 43316
rect 65828 43260 65838 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 76738 42924 76748 42980
rect 76804 42924 77420 42980
rect 77476 42924 77486 42980
rect 57922 42812 57932 42868
rect 57988 42812 58940 42868
rect 58996 42812 60396 42868
rect 60452 42812 60462 42868
rect 62738 42812 62748 42868
rect 62804 42812 63868 42868
rect 63924 42812 63934 42868
rect 67218 42812 67228 42868
rect 67284 42812 68572 42868
rect 68628 42812 69356 42868
rect 69412 42812 69422 42868
rect 80546 42812 80556 42868
rect 80612 42812 90076 42868
rect 90132 42812 90142 42868
rect 94322 42812 94332 42868
rect 94388 42812 94556 42868
rect 94612 42812 95564 42868
rect 95620 42812 96124 42868
rect 96180 42812 96190 42868
rect 75730 42700 75740 42756
rect 75796 42700 77756 42756
rect 77812 42700 77980 42756
rect 78036 42700 78046 42756
rect 86146 42700 86156 42756
rect 86212 42700 86716 42756
rect 86772 42700 89740 42756
rect 89796 42700 89806 42756
rect 92306 42700 92316 42756
rect 92372 42700 93212 42756
rect 93268 42700 93278 42756
rect 78530 42588 78540 42644
rect 78596 42588 79548 42644
rect 79604 42588 79614 42644
rect 84130 42588 84140 42644
rect 84196 42588 85260 42644
rect 85316 42588 86380 42644
rect 86436 42588 86446 42644
rect 73266 42476 73276 42532
rect 73332 42476 75180 42532
rect 75236 42476 76188 42532
rect 76244 42476 76254 42532
rect 86594 42476 86604 42532
rect 86660 42476 88284 42532
rect 88340 42476 89292 42532
rect 89348 42476 89358 42532
rect 92418 42476 92428 42532
rect 92484 42476 95004 42532
rect 95060 42476 95340 42532
rect 95396 42476 95406 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 78932 42140 88732 42196
rect 88788 42140 89964 42196
rect 90020 42140 92988 42196
rect 93044 42140 94052 42196
rect 78932 42084 78988 42140
rect 52658 42028 52668 42084
rect 52724 42028 54124 42084
rect 54180 42028 54684 42084
rect 54740 42028 54750 42084
rect 64652 42028 65772 42084
rect 65828 42028 65838 42084
rect 77746 42028 77756 42084
rect 77812 42028 78988 42084
rect 83906 42028 83916 42084
rect 83972 42028 84700 42084
rect 84756 42028 88508 42084
rect 88564 42028 92652 42084
rect 92708 42028 92718 42084
rect 56466 41916 56476 41972
rect 56532 41916 56542 41972
rect 57026 41916 57036 41972
rect 57092 41916 57596 41972
rect 57652 41916 60732 41972
rect 60788 41916 61292 41972
rect 61348 41916 61852 41972
rect 61908 41916 61918 41972
rect 56476 41860 56532 41916
rect 64652 41860 64708 42028
rect 93996 41972 94052 42140
rect 71698 41916 71708 41972
rect 71764 41916 73276 41972
rect 73332 41916 73342 41972
rect 93996 41916 95228 41972
rect 95284 41916 98028 41972
rect 98084 41916 98094 41972
rect 71708 41860 71764 41916
rect 51762 41804 51772 41860
rect 51828 41804 52444 41860
rect 52500 41804 53452 41860
rect 53508 41804 53518 41860
rect 56476 41804 56924 41860
rect 56980 41804 56990 41860
rect 60162 41804 60172 41860
rect 60228 41804 63420 41860
rect 63476 41804 63486 41860
rect 64642 41804 64652 41860
rect 64708 41804 64718 41860
rect 68674 41804 68684 41860
rect 68740 41804 69244 41860
rect 69300 41804 70476 41860
rect 70532 41804 70542 41860
rect 70802 41804 70812 41860
rect 70868 41804 71764 41860
rect 77410 41804 77420 41860
rect 77476 41804 78204 41860
rect 78260 41804 78270 41860
rect 92642 41804 92652 41860
rect 92708 41804 94332 41860
rect 94388 41804 95676 41860
rect 95732 41804 95742 41860
rect 61730 41692 61740 41748
rect 61796 41692 62412 41748
rect 62468 41692 64316 41748
rect 64372 41692 64382 41748
rect 75282 41692 75292 41748
rect 75348 41692 77308 41748
rect 77364 41692 77374 41748
rect 94882 41692 94892 41748
rect 94948 41692 96012 41748
rect 96068 41692 96078 41748
rect 70690 41580 70700 41636
rect 70756 41580 72268 41636
rect 72324 41580 72334 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 64306 41468 64316 41524
rect 64372 41468 65436 41524
rect 65492 41468 65502 41524
rect 55132 41356 56924 41412
rect 56980 41356 72268 41412
rect 72324 41356 74060 41412
rect 74116 41356 74126 41412
rect 89730 41356 89740 41412
rect 89796 41356 90300 41412
rect 90356 41356 90366 41412
rect 55132 41300 55188 41356
rect 52546 41244 52556 41300
rect 52612 41244 54236 41300
rect 54292 41244 55132 41300
rect 55188 41244 55198 41300
rect 62178 41244 62188 41300
rect 62244 41244 64204 41300
rect 64260 41244 64270 41300
rect 64418 41244 64428 41300
rect 64484 41244 65548 41300
rect 65604 41244 69468 41300
rect 69524 41244 70364 41300
rect 70420 41244 70924 41300
rect 70980 41244 70990 41300
rect 75842 41244 75852 41300
rect 75908 41244 76524 41300
rect 76580 41244 80556 41300
rect 80612 41244 80622 41300
rect 89842 41244 89852 41300
rect 89908 41244 90412 41300
rect 90468 41244 90478 41300
rect 93538 41244 93548 41300
rect 93604 41244 95340 41300
rect 95396 41244 95406 41300
rect 50754 41132 50764 41188
rect 50820 41132 53116 41188
rect 53172 41132 53182 41188
rect 57698 41132 57708 41188
rect 57764 41132 58604 41188
rect 58660 41132 58670 41188
rect 63074 41132 63084 41188
rect 63140 41132 64988 41188
rect 65044 41132 65996 41188
rect 66052 41132 66444 41188
rect 66500 41132 66510 41188
rect 67666 41132 67676 41188
rect 67732 41132 69916 41188
rect 69972 41132 69982 41188
rect 71250 41132 71260 41188
rect 71316 41132 71820 41188
rect 71876 41132 72716 41188
rect 72772 41132 73948 41188
rect 74610 41132 74620 41188
rect 74676 41132 75292 41188
rect 75348 41132 75358 41188
rect 89618 41132 89628 41188
rect 89684 41132 90748 41188
rect 90804 41132 90814 41188
rect 91298 41132 91308 41188
rect 91364 41132 97356 41188
rect 97412 41132 97580 41188
rect 97636 41132 97646 41188
rect 65548 41076 65604 41132
rect 72268 41076 72324 41132
rect 49522 41020 49532 41076
rect 49588 41020 51436 41076
rect 51492 41020 51502 41076
rect 52322 41020 52332 41076
rect 52388 41020 54684 41076
rect 54740 41020 62748 41076
rect 62804 41020 62814 41076
rect 65538 41020 65548 41076
rect 65604 41020 65614 41076
rect 72258 41020 72268 41076
rect 72324 41020 72334 41076
rect 73892 40964 73948 41132
rect 74722 41020 74732 41076
rect 74788 41020 77308 41076
rect 77364 41020 77374 41076
rect 81554 41020 81564 41076
rect 81620 41020 81788 41076
rect 81844 41020 82684 41076
rect 82740 41020 82750 41076
rect 83234 41020 83244 41076
rect 83300 41020 84252 41076
rect 84308 41020 84318 41076
rect 92418 41020 92428 41076
rect 92484 41020 96796 41076
rect 96852 41020 96862 41076
rect 58146 40908 58156 40964
rect 58212 40908 59500 40964
rect 59556 40908 59566 40964
rect 69906 40908 69916 40964
rect 69972 40908 70812 40964
rect 70868 40908 70878 40964
rect 73892 40908 75292 40964
rect 75348 40908 76300 40964
rect 76356 40908 76366 40964
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 62178 40572 62188 40628
rect 62244 40572 63084 40628
rect 63140 40572 63150 40628
rect 88834 40572 88844 40628
rect 88900 40572 89292 40628
rect 89348 40572 89358 40628
rect 96338 40572 96348 40628
rect 96404 40572 97468 40628
rect 97524 40572 97534 40628
rect 62738 40460 62748 40516
rect 62804 40460 63532 40516
rect 63588 40460 63598 40516
rect 63970 40460 63980 40516
rect 64036 40460 65212 40516
rect 65268 40460 65278 40516
rect 73938 40460 73948 40516
rect 74004 40460 75516 40516
rect 75572 40460 77756 40516
rect 77812 40460 78204 40516
rect 78260 40460 78270 40516
rect 93650 40460 93660 40516
rect 93716 40460 93996 40516
rect 94052 40460 96124 40516
rect 96180 40460 96908 40516
rect 96964 40460 96974 40516
rect 55570 40348 55580 40404
rect 55636 40348 56028 40404
rect 56084 40348 57036 40404
rect 57092 40348 57102 40404
rect 58930 40348 58940 40404
rect 58996 40348 61292 40404
rect 61348 40348 61358 40404
rect 72034 40348 72044 40404
rect 72100 40348 77196 40404
rect 77252 40348 77262 40404
rect 80434 40348 80444 40404
rect 80500 40348 81228 40404
rect 81284 40348 83916 40404
rect 83972 40348 83982 40404
rect 82450 40236 82460 40292
rect 82516 40236 83804 40292
rect 83860 40236 83870 40292
rect 84914 40236 84924 40292
rect 84980 40236 85820 40292
rect 85876 40236 88172 40292
rect 88228 40236 88238 40292
rect 82674 40124 82684 40180
rect 82740 40124 84140 40180
rect 84196 40124 84206 40180
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 70242 39676 70252 39732
rect 70308 39676 70700 39732
rect 70756 39676 71260 39732
rect 71316 39676 71326 39732
rect 73826 39676 73836 39732
rect 73892 39676 74844 39732
rect 74900 39676 75180 39732
rect 75236 39676 75246 39732
rect 81330 39676 81340 39732
rect 81396 39676 82908 39732
rect 82964 39676 82974 39732
rect 83794 39676 83804 39732
rect 83860 39676 87948 39732
rect 88004 39676 90636 39732
rect 90692 39676 90702 39732
rect 94882 39676 94892 39732
rect 94948 39676 95340 39732
rect 95396 39676 98252 39732
rect 98308 39676 98318 39732
rect 60722 39564 60732 39620
rect 60788 39564 61740 39620
rect 61796 39564 62300 39620
rect 62356 39564 62366 39620
rect 75394 39564 75404 39620
rect 75460 39564 76412 39620
rect 76468 39564 77308 39620
rect 77364 39564 77374 39620
rect 82338 39564 82348 39620
rect 82404 39564 83244 39620
rect 83300 39564 83310 39620
rect 51426 39452 51436 39508
rect 51492 39452 52332 39508
rect 52388 39452 53676 39508
rect 53732 39452 53742 39508
rect 14242 39340 14252 39396
rect 14308 39340 50540 39396
rect 50596 39340 51100 39396
rect 51156 39340 51166 39396
rect 60274 39340 60284 39396
rect 60340 39340 62188 39396
rect 62514 39340 62524 39396
rect 62580 39340 63756 39396
rect 63812 39340 63822 39396
rect 62132 39284 62188 39340
rect 62132 39228 63196 39284
rect 63252 39228 63262 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 59938 39004 59948 39060
rect 60004 39004 62188 39060
rect 62244 39004 62254 39060
rect 68562 39004 68572 39060
rect 68628 39004 69692 39060
rect 69748 39004 69758 39060
rect 70690 39004 70700 39060
rect 70756 39004 71372 39060
rect 71428 39004 71932 39060
rect 71988 39004 78988 39060
rect 81442 39004 81452 39060
rect 81508 39004 82572 39060
rect 82628 39004 84476 39060
rect 84532 39004 85148 39060
rect 85204 39004 85820 39060
rect 85876 39004 85886 39060
rect 54562 38892 54572 38948
rect 54628 38892 55468 38948
rect 55524 38892 55534 38948
rect 62850 38892 62860 38948
rect 62916 38892 63980 38948
rect 64036 38892 64046 38948
rect 74834 38892 74844 38948
rect 74900 38892 76188 38948
rect 76244 38892 76254 38948
rect 78932 38836 78988 39004
rect 80098 38892 80108 38948
rect 80164 38892 81116 38948
rect 81172 38892 81182 38948
rect 90178 38892 90188 38948
rect 90244 38892 91532 38948
rect 91588 38892 91598 38948
rect 52892 38780 53452 38836
rect 53508 38780 53788 38836
rect 53844 38780 53854 38836
rect 63410 38780 63420 38836
rect 63476 38780 64204 38836
rect 64260 38780 64270 38836
rect 74946 38780 74956 38836
rect 75012 38780 77532 38836
rect 77588 38780 77598 38836
rect 78932 38780 82460 38836
rect 82516 38780 82526 38836
rect 91186 38780 91196 38836
rect 91252 38780 93100 38836
rect 93156 38780 94220 38836
rect 94276 38780 94286 38836
rect 96450 38780 96460 38836
rect 96516 38780 97468 38836
rect 97524 38780 97534 38836
rect 52892 38724 52948 38780
rect 52882 38668 52892 38724
rect 52948 38668 52958 38724
rect 61506 38668 61516 38724
rect 61572 38668 62524 38724
rect 62580 38668 62590 38724
rect 63186 38668 63196 38724
rect 63252 38668 65660 38724
rect 65716 38668 65726 38724
rect 68226 38668 68236 38724
rect 68292 38668 69804 38724
rect 69860 38668 69870 38724
rect 75618 38668 75628 38724
rect 75684 38668 78316 38724
rect 78372 38668 79324 38724
rect 79380 38668 79390 38724
rect 95778 38668 95788 38724
rect 95844 38668 97020 38724
rect 97076 38668 98028 38724
rect 98084 38668 98094 38724
rect 93874 38556 93884 38612
rect 93940 38556 94332 38612
rect 94388 38556 95452 38612
rect 95508 38556 96236 38612
rect 96292 38556 98140 38612
rect 98196 38556 98206 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 52658 38108 52668 38164
rect 52724 38108 53452 38164
rect 53508 38108 53518 38164
rect 61058 38108 61068 38164
rect 61124 38108 61516 38164
rect 61572 38108 63084 38164
rect 63140 38108 63150 38164
rect 68338 38108 68348 38164
rect 68404 38108 69244 38164
rect 69300 38108 69310 38164
rect 77746 38108 77756 38164
rect 77812 38108 78988 38164
rect 79044 38108 79054 38164
rect 83234 38108 83244 38164
rect 83300 38108 83580 38164
rect 83636 38108 84252 38164
rect 84308 38108 84318 38164
rect 61282 37996 61292 38052
rect 61348 37996 62188 38052
rect 62244 37996 64540 38052
rect 64596 37996 65324 38052
rect 65380 37996 65390 38052
rect 67554 37996 67564 38052
rect 67620 37996 69580 38052
rect 69636 37996 69646 38052
rect 75842 37996 75852 38052
rect 75908 37996 76524 38052
rect 76580 37996 76590 38052
rect 77858 37996 77868 38052
rect 77924 37996 78540 38052
rect 78596 37996 79996 38052
rect 80052 37996 80062 38052
rect 89506 37996 89516 38052
rect 89572 37996 91644 38052
rect 91700 37996 91710 38052
rect 66546 37884 66556 37940
rect 66612 37884 67228 37940
rect 67284 37884 67294 37940
rect 75954 37884 75964 37940
rect 76020 37884 77084 37940
rect 77140 37884 77150 37940
rect 94098 37884 94108 37940
rect 94164 37884 95452 37940
rect 95508 37884 95518 37940
rect 55682 37772 55692 37828
rect 55748 37772 57260 37828
rect 57316 37772 58156 37828
rect 58212 37772 61516 37828
rect 61572 37772 61582 37828
rect 79986 37772 79996 37828
rect 80052 37772 88508 37828
rect 88564 37772 90972 37828
rect 91028 37772 91038 37828
rect 57362 37660 57372 37716
rect 57428 37660 58044 37716
rect 58100 37660 58716 37716
rect 58772 37660 59388 37716
rect 59444 37660 59724 37716
rect 59780 37660 68348 37716
rect 68404 37660 68414 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 0 37492 800 37520
rect 0 37436 1820 37492
rect 1876 37436 1886 37492
rect 58818 37436 58828 37492
rect 58884 37436 59836 37492
rect 59892 37436 61180 37492
rect 61236 37436 61246 37492
rect 0 37408 800 37436
rect 49186 37324 49196 37380
rect 49252 37324 50316 37380
rect 50372 37324 50382 37380
rect 64418 37324 64428 37380
rect 64484 37324 64988 37380
rect 65044 37324 65212 37380
rect 65268 37324 75852 37380
rect 75908 37324 77868 37380
rect 77924 37324 77934 37380
rect 89394 37324 89404 37380
rect 89460 37324 91420 37380
rect 91476 37324 91486 37380
rect 91970 37324 91980 37380
rect 92036 37324 93100 37380
rect 93156 37324 93166 37380
rect 56466 37212 56476 37268
rect 56532 37212 57708 37268
rect 57764 37212 57774 37268
rect 66770 37212 66780 37268
rect 66836 37212 70140 37268
rect 70196 37212 70206 37268
rect 82226 37212 82236 37268
rect 82292 37212 82908 37268
rect 82964 37212 82974 37268
rect 95554 37212 95564 37268
rect 95620 37212 96012 37268
rect 96068 37212 97580 37268
rect 97636 37212 97646 37268
rect 51426 37100 51436 37156
rect 51492 37100 52444 37156
rect 52500 37100 52510 37156
rect 83794 37100 83804 37156
rect 83860 37100 84588 37156
rect 84644 37100 84654 37156
rect 89282 37100 89292 37156
rect 89348 37100 90300 37156
rect 90356 37100 90366 37156
rect 61506 36988 61516 37044
rect 61572 36988 61964 37044
rect 62020 36988 62030 37044
rect 91634 36988 91644 37044
rect 91700 36988 92764 37044
rect 92820 36988 92830 37044
rect 73378 36876 73388 36932
rect 73444 36876 74060 36932
rect 74116 36876 74620 36932
rect 74676 36876 75404 36932
rect 75460 36876 75470 36932
rect 76402 36876 76412 36932
rect 76468 36876 77196 36932
rect 77252 36876 77532 36932
rect 77588 36876 77598 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 70578 36764 70588 36820
rect 70644 36764 71148 36820
rect 71204 36764 71708 36820
rect 71764 36764 81788 36820
rect 81844 36764 81854 36820
rect 48962 36652 48972 36708
rect 49028 36652 51100 36708
rect 51156 36652 51166 36708
rect 93762 36652 93772 36708
rect 93828 36652 95228 36708
rect 95284 36652 95294 36708
rect 54338 36540 54348 36596
rect 54404 36540 55580 36596
rect 55636 36540 55646 36596
rect 76066 36540 76076 36596
rect 76132 36540 77420 36596
rect 77476 36540 77644 36596
rect 77700 36540 77710 36596
rect 86706 36540 86716 36596
rect 86772 36540 87052 36596
rect 87108 36540 88172 36596
rect 88228 36540 88732 36596
rect 88788 36540 88798 36596
rect 90962 36540 90972 36596
rect 91028 36540 93212 36596
rect 93268 36540 95452 36596
rect 95508 36540 95788 36596
rect 95844 36540 97132 36596
rect 97188 36540 97198 36596
rect 52210 36428 52220 36484
rect 52276 36428 52780 36484
rect 52836 36428 53340 36484
rect 53396 36428 54124 36484
rect 54180 36428 54190 36484
rect 74610 36428 74620 36484
rect 74676 36428 74956 36484
rect 75012 36428 84924 36484
rect 84980 36428 84990 36484
rect 93762 36428 93772 36484
rect 93828 36428 95340 36484
rect 95396 36428 95406 36484
rect 52098 36316 52108 36372
rect 52164 36316 53676 36372
rect 53732 36316 53742 36372
rect 68338 36316 68348 36372
rect 68404 36316 69468 36372
rect 69524 36316 69534 36372
rect 70354 36316 70364 36372
rect 70420 36316 70812 36372
rect 70868 36316 71596 36372
rect 71652 36316 71662 36372
rect 74946 36204 74956 36260
rect 75012 36204 76412 36260
rect 76468 36204 76478 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 62738 35980 62748 36036
rect 62804 35980 63756 36036
rect 63812 35980 64316 36036
rect 64372 35980 64382 36036
rect 54114 35868 54124 35924
rect 54180 35868 55244 35924
rect 55300 35868 74284 35924
rect 74340 35868 74732 35924
rect 74788 35868 75292 35924
rect 75348 35868 75358 35924
rect 81218 35868 81228 35924
rect 81284 35868 81788 35924
rect 81844 35868 81854 35924
rect 58034 35756 58044 35812
rect 58100 35756 58604 35812
rect 58660 35756 61068 35812
rect 61124 35756 61134 35812
rect 74386 35756 74396 35812
rect 74452 35756 76524 35812
rect 76580 35756 76590 35812
rect 84914 35756 84924 35812
rect 84980 35756 86156 35812
rect 86212 35756 87948 35812
rect 88004 35756 88508 35812
rect 88564 35756 89964 35812
rect 90020 35756 90030 35812
rect 52882 35644 52892 35700
rect 52948 35644 53564 35700
rect 53620 35644 54460 35700
rect 54516 35644 54526 35700
rect 60274 35644 60284 35700
rect 60340 35644 63084 35700
rect 63140 35644 63150 35700
rect 61730 35532 61740 35588
rect 61796 35532 66668 35588
rect 66724 35532 67228 35588
rect 67284 35532 67294 35588
rect 51314 35420 51324 35476
rect 51380 35420 53564 35476
rect 53620 35420 53630 35476
rect 57474 35420 57484 35476
rect 57540 35420 58156 35476
rect 58212 35420 58716 35476
rect 58772 35420 58782 35476
rect 52658 35308 52668 35364
rect 52724 35308 53900 35364
rect 53956 35308 53966 35364
rect 81778 35308 81788 35364
rect 81844 35308 82292 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 82236 35252 82292 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 82236 35196 82908 35252
rect 82964 35196 82974 35252
rect 92866 35196 92876 35252
rect 92932 35196 96124 35252
rect 96180 35196 96190 35252
rect 56690 34972 56700 35028
rect 56756 34972 57372 35028
rect 57428 34972 57438 35028
rect 60610 34972 60620 35028
rect 60676 34972 62188 35028
rect 62244 34972 62254 35028
rect 62514 34972 62524 35028
rect 62580 34972 63644 35028
rect 63700 34972 66108 35028
rect 66164 34972 66668 35028
rect 66724 34972 72380 35028
rect 72436 34972 73500 35028
rect 73556 34972 73566 35028
rect 75506 34972 75516 35028
rect 75572 34972 76524 35028
rect 76580 34972 77084 35028
rect 77140 34972 77150 35028
rect 49858 34860 49868 34916
rect 49924 34860 53676 34916
rect 53732 34860 53742 34916
rect 63858 34860 63868 34916
rect 63924 34860 65324 34916
rect 65380 34860 65390 34916
rect 68226 34860 68236 34916
rect 68292 34860 68572 34916
rect 68628 34860 69692 34916
rect 69748 34860 69758 34916
rect 72146 34860 72156 34916
rect 72212 34860 72604 34916
rect 72660 34860 72670 34916
rect 73714 34860 73724 34916
rect 73780 34860 77308 34916
rect 77364 34860 77756 34916
rect 77812 34860 77822 34916
rect 82114 34860 82124 34916
rect 82180 34860 82684 34916
rect 82740 34860 82750 34916
rect 84242 34860 84252 34916
rect 84308 34860 85596 34916
rect 85652 34860 85662 34916
rect 89506 34860 89516 34916
rect 89572 34860 91644 34916
rect 91700 34860 91710 34916
rect 52994 34748 53004 34804
rect 53060 34748 54012 34804
rect 54068 34748 54684 34804
rect 54740 34748 55692 34804
rect 55748 34748 55758 34804
rect 81666 34748 81676 34804
rect 81732 34748 83244 34804
rect 83300 34748 83310 34804
rect 84466 34748 84476 34804
rect 84532 34748 86044 34804
rect 86100 34748 86110 34804
rect 59938 34636 59948 34692
rect 60004 34636 68460 34692
rect 68516 34636 69356 34692
rect 69412 34636 72044 34692
rect 72100 34636 72110 34692
rect 88050 34636 88060 34692
rect 88116 34636 88620 34692
rect 88676 34636 88686 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 85138 34412 85148 34468
rect 85204 34412 85932 34468
rect 85988 34412 87500 34468
rect 87556 34412 87566 34468
rect 90692 34412 90972 34468
rect 91028 34412 93660 34468
rect 93716 34412 93996 34468
rect 94052 34412 94062 34468
rect 90692 34356 90748 34412
rect 62178 34300 62188 34356
rect 62244 34300 63308 34356
rect 63364 34300 64540 34356
rect 64596 34300 65884 34356
rect 65940 34300 65950 34356
rect 71138 34300 71148 34356
rect 71204 34300 73500 34356
rect 73556 34300 73566 34356
rect 77522 34300 77532 34356
rect 77588 34300 89852 34356
rect 89908 34300 90748 34356
rect 94322 34300 94332 34356
rect 94388 34300 95228 34356
rect 95284 34300 95294 34356
rect 96114 34300 96124 34356
rect 96180 34300 97132 34356
rect 97188 34300 97468 34356
rect 97524 34300 97534 34356
rect 56690 34188 56700 34244
rect 56756 34188 56766 34244
rect 64978 34188 64988 34244
rect 65044 34188 65772 34244
rect 65828 34188 65838 34244
rect 79874 34188 79884 34244
rect 79940 34188 82348 34244
rect 82404 34188 82414 34244
rect 86482 34188 86492 34244
rect 86548 34188 87612 34244
rect 87668 34188 87678 34244
rect 91970 34188 91980 34244
rect 92036 34188 93100 34244
rect 93156 34188 93166 34244
rect 56700 34132 56756 34188
rect 53890 34076 53900 34132
rect 53956 34076 54460 34132
rect 54516 34076 58268 34132
rect 58324 34076 60284 34132
rect 60340 34076 60732 34132
rect 60788 34076 60956 34132
rect 61012 34076 61022 34132
rect 72594 34076 72604 34132
rect 72660 34076 73836 34132
rect 73892 34076 73902 34132
rect 78754 34076 78764 34132
rect 78820 34076 82460 34132
rect 82516 34076 82526 34132
rect 85810 34076 85820 34132
rect 85876 34076 86604 34132
rect 86660 34076 86940 34132
rect 86996 34076 88396 34132
rect 88452 34076 89180 34132
rect 89236 34076 89246 34132
rect 89394 34076 89404 34132
rect 89460 34076 92428 34132
rect 92484 34076 92494 34132
rect 95554 34076 95564 34132
rect 95620 34076 97244 34132
rect 97300 34076 97310 34132
rect 56690 33964 56700 34020
rect 56756 33964 57932 34020
rect 57988 33964 58380 34020
rect 58436 33964 58446 34020
rect 61954 33964 61964 34020
rect 62020 33964 63868 34020
rect 63924 33964 63934 34020
rect 90738 33964 90748 34020
rect 90804 33964 92204 34020
rect 92260 33964 92270 34020
rect 83906 33852 83916 33908
rect 83972 33852 87276 33908
rect 87332 33852 87342 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 77868 33628 79436 33684
rect 79492 33628 79502 33684
rect 81106 33628 81116 33684
rect 81172 33628 82124 33684
rect 82180 33628 82190 33684
rect 86706 33628 86716 33684
rect 86772 33628 87836 33684
rect 87892 33628 87902 33684
rect 89506 33628 89516 33684
rect 89572 33628 90188 33684
rect 90244 33628 90254 33684
rect 91634 33628 91644 33684
rect 91700 33628 92764 33684
rect 92820 33628 92830 33684
rect 77868 33572 77924 33628
rect 77858 33516 77868 33572
rect 77924 33516 77934 33572
rect 93986 33516 93996 33572
rect 94052 33516 95788 33572
rect 95844 33516 95854 33572
rect 53106 33404 53116 33460
rect 53172 33404 53788 33460
rect 53844 33404 55468 33460
rect 55412 33236 55468 33404
rect 57362 33292 57372 33348
rect 57428 33292 58380 33348
rect 58436 33292 58446 33348
rect 59154 33292 59164 33348
rect 59220 33292 59724 33348
rect 59780 33292 59790 33348
rect 64978 33292 64988 33348
rect 65044 33292 65772 33348
rect 65828 33292 66332 33348
rect 66388 33292 68684 33348
rect 68740 33292 69692 33348
rect 69748 33292 70812 33348
rect 70868 33292 70878 33348
rect 73714 33292 73724 33348
rect 73780 33292 74732 33348
rect 74788 33292 74798 33348
rect 76290 33292 76300 33348
rect 76356 33292 77532 33348
rect 77588 33292 77598 33348
rect 80658 33292 80668 33348
rect 80724 33292 82796 33348
rect 82852 33292 82862 33348
rect 92418 33292 92428 33348
rect 92484 33292 94444 33348
rect 94500 33292 94510 33348
rect 59164 33236 59220 33292
rect 55412 33180 56476 33236
rect 56532 33180 57036 33236
rect 57092 33180 59220 33236
rect 60610 33180 60620 33236
rect 60676 33180 61740 33236
rect 61796 33180 61806 33236
rect 70354 33180 70364 33236
rect 70420 33180 71372 33236
rect 71428 33180 74284 33236
rect 74340 33180 85596 33236
rect 85652 33180 85662 33236
rect 55906 33068 55916 33124
rect 55972 33068 58044 33124
rect 58100 33068 58110 33124
rect 70242 33068 70252 33124
rect 70308 33068 73052 33124
rect 73108 33068 73836 33124
rect 73892 33068 73902 33124
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 57810 32732 57820 32788
rect 57876 32732 58940 32788
rect 58996 32732 59724 32788
rect 59780 32732 59790 32788
rect 60386 32732 60396 32788
rect 60452 32732 61740 32788
rect 61796 32732 61806 32788
rect 72594 32732 72604 32788
rect 72660 32732 73836 32788
rect 73892 32732 74284 32788
rect 74340 32732 75516 32788
rect 75572 32732 75582 32788
rect 76738 32732 76748 32788
rect 76804 32732 77308 32788
rect 77364 32732 77374 32788
rect 78978 32732 78988 32788
rect 79044 32732 81340 32788
rect 81396 32732 81406 32788
rect 82898 32732 82908 32788
rect 82964 32732 83692 32788
rect 83748 32732 84364 32788
rect 84420 32732 86044 32788
rect 86100 32732 88172 32788
rect 88228 32732 88238 32788
rect 94658 32732 94668 32788
rect 94724 32732 96236 32788
rect 96292 32732 96302 32788
rect 59724 32676 59780 32732
rect 59724 32620 61404 32676
rect 61460 32620 62636 32676
rect 62692 32620 62702 32676
rect 76178 32620 76188 32676
rect 76244 32620 77868 32676
rect 77924 32620 77934 32676
rect 85586 32620 85596 32676
rect 85652 32620 87388 32676
rect 87444 32620 90748 32676
rect 90692 32564 90748 32620
rect 54786 32508 54796 32564
rect 54852 32508 55468 32564
rect 55524 32508 55534 32564
rect 55794 32508 55804 32564
rect 55860 32508 57372 32564
rect 57428 32508 57438 32564
rect 70914 32508 70924 32564
rect 70980 32508 73276 32564
rect 73332 32508 73342 32564
rect 90692 32508 90972 32564
rect 91028 32508 91532 32564
rect 91588 32508 91598 32564
rect 67666 32396 67676 32452
rect 67732 32396 68572 32452
rect 68628 32396 69580 32452
rect 69636 32396 69646 32452
rect 68002 32284 68012 32340
rect 68068 32284 69244 32340
rect 69300 32284 69310 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 89282 31836 89292 31892
rect 89348 31836 90748 31892
rect 90804 31836 90814 31892
rect 67442 31724 67452 31780
rect 67508 31724 69356 31780
rect 69412 31724 69422 31780
rect 66434 31612 66444 31668
rect 66500 31612 67676 31668
rect 67732 31612 67742 31668
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 82338 30940 82348 30996
rect 82404 30940 83132 30996
rect 83188 30940 83198 30996
rect 84578 30828 84588 30884
rect 84644 30828 86044 30884
rect 86100 30828 87052 30884
rect 87108 30828 87118 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 83682 29484 83692 29540
rect 83748 29484 85148 29540
rect 85204 29484 85214 29540
rect 83234 29372 83244 29428
rect 83300 29372 85372 29428
rect 85428 29372 85438 29428
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 76962 25228 76972 25284
rect 77028 25228 94892 25284
rect 94948 25228 94958 25284
rect 95218 25228 95228 25284
rect 95284 25228 95788 25284
rect 95844 25228 95854 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 95788 25060 95844 25228
rect 99200 25060 100000 25088
rect 95788 25004 100000 25060
rect 99200 24976 100000 25004
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 2146 12684 2156 12740
rect 2212 12684 73388 12740
rect 73444 12684 73454 12740
rect 0 12516 800 12544
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 0 12460 1820 12516
rect 1876 12460 1886 12516
rect 0 12432 800 12460
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 43698 3388 43708 3444
rect 43764 3388 44268 3444
rect 44324 3388 44940 3444
rect 44996 3388 45006 3444
rect 56130 3388 56140 3444
rect 56196 3388 56700 3444
rect 56756 3388 56766 3444
rect 67778 3388 67788 3444
rect 67844 3388 68796 3444
rect 68852 3388 68862 3444
rect 93426 3388 93436 3444
rect 93492 3388 93996 3444
rect 94052 3388 94062 3444
rect 6962 3276 6972 3332
rect 7028 3276 14252 3332
rect 14308 3276 14318 3332
rect 19394 3276 19404 3332
rect 19460 3276 54348 3332
rect 54404 3276 54414 3332
rect 69122 3276 69132 3332
rect 69188 3276 89628 3332
rect 89684 3276 89694 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 57026 2940 57036 2996
rect 57092 2940 82460 2996
rect 82516 2940 82526 2996
rect 31826 2828 31836 2884
rect 31892 2828 57372 2884
rect 57428 2828 57438 2884
rect 77522 2828 77532 2884
rect 77588 2828 93660 2884
rect 93716 2828 93726 2884
rect 45266 2716 45276 2772
rect 45332 2716 69020 2772
rect 69076 2716 69086 2772
<< via3 >>
rect 4476 96404 4532 96460
rect 4580 96404 4636 96460
rect 4684 96404 4740 96460
rect 35196 96404 35252 96460
rect 35300 96404 35356 96460
rect 35404 96404 35460 96460
rect 65916 96404 65972 96460
rect 66020 96404 66076 96460
rect 66124 96404 66180 96460
rect 96636 96404 96692 96460
rect 96740 96404 96796 96460
rect 96844 96404 96900 96460
rect 19836 95620 19892 95676
rect 19940 95620 19996 95676
rect 20044 95620 20100 95676
rect 50556 95620 50612 95676
rect 50660 95620 50716 95676
rect 50764 95620 50820 95676
rect 81276 95620 81332 95676
rect 81380 95620 81436 95676
rect 81484 95620 81540 95676
rect 4476 94836 4532 94892
rect 4580 94836 4636 94892
rect 4684 94836 4740 94892
rect 35196 94836 35252 94892
rect 35300 94836 35356 94892
rect 35404 94836 35460 94892
rect 65916 94836 65972 94892
rect 66020 94836 66076 94892
rect 66124 94836 66180 94892
rect 96636 94836 96692 94892
rect 96740 94836 96796 94892
rect 96844 94836 96900 94892
rect 19836 94052 19892 94108
rect 19940 94052 19996 94108
rect 20044 94052 20100 94108
rect 50556 94052 50612 94108
rect 50660 94052 50716 94108
rect 50764 94052 50820 94108
rect 81276 94052 81332 94108
rect 81380 94052 81436 94108
rect 81484 94052 81540 94108
rect 4476 93268 4532 93324
rect 4580 93268 4636 93324
rect 4684 93268 4740 93324
rect 35196 93268 35252 93324
rect 35300 93268 35356 93324
rect 35404 93268 35460 93324
rect 65916 93268 65972 93324
rect 66020 93268 66076 93324
rect 66124 93268 66180 93324
rect 96636 93268 96692 93324
rect 96740 93268 96796 93324
rect 96844 93268 96900 93324
rect 19836 92484 19892 92540
rect 19940 92484 19996 92540
rect 20044 92484 20100 92540
rect 50556 92484 50612 92540
rect 50660 92484 50716 92540
rect 50764 92484 50820 92540
rect 81276 92484 81332 92540
rect 81380 92484 81436 92540
rect 81484 92484 81540 92540
rect 4476 91700 4532 91756
rect 4580 91700 4636 91756
rect 4684 91700 4740 91756
rect 35196 91700 35252 91756
rect 35300 91700 35356 91756
rect 35404 91700 35460 91756
rect 65916 91700 65972 91756
rect 66020 91700 66076 91756
rect 66124 91700 66180 91756
rect 96636 91700 96692 91756
rect 96740 91700 96796 91756
rect 96844 91700 96900 91756
rect 19836 90916 19892 90972
rect 19940 90916 19996 90972
rect 20044 90916 20100 90972
rect 50556 90916 50612 90972
rect 50660 90916 50716 90972
rect 50764 90916 50820 90972
rect 81276 90916 81332 90972
rect 81380 90916 81436 90972
rect 81484 90916 81540 90972
rect 4476 90132 4532 90188
rect 4580 90132 4636 90188
rect 4684 90132 4740 90188
rect 35196 90132 35252 90188
rect 35300 90132 35356 90188
rect 35404 90132 35460 90188
rect 65916 90132 65972 90188
rect 66020 90132 66076 90188
rect 66124 90132 66180 90188
rect 96636 90132 96692 90188
rect 96740 90132 96796 90188
rect 96844 90132 96900 90188
rect 19836 89348 19892 89404
rect 19940 89348 19996 89404
rect 20044 89348 20100 89404
rect 50556 89348 50612 89404
rect 50660 89348 50716 89404
rect 50764 89348 50820 89404
rect 81276 89348 81332 89404
rect 81380 89348 81436 89404
rect 81484 89348 81540 89404
rect 4476 88564 4532 88620
rect 4580 88564 4636 88620
rect 4684 88564 4740 88620
rect 35196 88564 35252 88620
rect 35300 88564 35356 88620
rect 35404 88564 35460 88620
rect 65916 88564 65972 88620
rect 66020 88564 66076 88620
rect 66124 88564 66180 88620
rect 96636 88564 96692 88620
rect 96740 88564 96796 88620
rect 96844 88564 96900 88620
rect 19836 87780 19892 87836
rect 19940 87780 19996 87836
rect 20044 87780 20100 87836
rect 50556 87780 50612 87836
rect 50660 87780 50716 87836
rect 50764 87780 50820 87836
rect 81276 87780 81332 87836
rect 81380 87780 81436 87836
rect 81484 87780 81540 87836
rect 4476 86996 4532 87052
rect 4580 86996 4636 87052
rect 4684 86996 4740 87052
rect 35196 86996 35252 87052
rect 35300 86996 35356 87052
rect 35404 86996 35460 87052
rect 65916 86996 65972 87052
rect 66020 86996 66076 87052
rect 66124 86996 66180 87052
rect 96636 86996 96692 87052
rect 96740 86996 96796 87052
rect 96844 86996 96900 87052
rect 19836 86212 19892 86268
rect 19940 86212 19996 86268
rect 20044 86212 20100 86268
rect 50556 86212 50612 86268
rect 50660 86212 50716 86268
rect 50764 86212 50820 86268
rect 81276 86212 81332 86268
rect 81380 86212 81436 86268
rect 81484 86212 81540 86268
rect 4476 85428 4532 85484
rect 4580 85428 4636 85484
rect 4684 85428 4740 85484
rect 35196 85428 35252 85484
rect 35300 85428 35356 85484
rect 35404 85428 35460 85484
rect 65916 85428 65972 85484
rect 66020 85428 66076 85484
rect 66124 85428 66180 85484
rect 96636 85428 96692 85484
rect 96740 85428 96796 85484
rect 96844 85428 96900 85484
rect 19836 84644 19892 84700
rect 19940 84644 19996 84700
rect 20044 84644 20100 84700
rect 50556 84644 50612 84700
rect 50660 84644 50716 84700
rect 50764 84644 50820 84700
rect 81276 84644 81332 84700
rect 81380 84644 81436 84700
rect 81484 84644 81540 84700
rect 4476 83860 4532 83916
rect 4580 83860 4636 83916
rect 4684 83860 4740 83916
rect 35196 83860 35252 83916
rect 35300 83860 35356 83916
rect 35404 83860 35460 83916
rect 65916 83860 65972 83916
rect 66020 83860 66076 83916
rect 66124 83860 66180 83916
rect 96636 83860 96692 83916
rect 96740 83860 96796 83916
rect 96844 83860 96900 83916
rect 19836 83076 19892 83132
rect 19940 83076 19996 83132
rect 20044 83076 20100 83132
rect 50556 83076 50612 83132
rect 50660 83076 50716 83132
rect 50764 83076 50820 83132
rect 81276 83076 81332 83132
rect 81380 83076 81436 83132
rect 81484 83076 81540 83132
rect 4476 82292 4532 82348
rect 4580 82292 4636 82348
rect 4684 82292 4740 82348
rect 35196 82292 35252 82348
rect 35300 82292 35356 82348
rect 35404 82292 35460 82348
rect 65916 82292 65972 82348
rect 66020 82292 66076 82348
rect 66124 82292 66180 82348
rect 96636 82292 96692 82348
rect 96740 82292 96796 82348
rect 96844 82292 96900 82348
rect 19836 81508 19892 81564
rect 19940 81508 19996 81564
rect 20044 81508 20100 81564
rect 50556 81508 50612 81564
rect 50660 81508 50716 81564
rect 50764 81508 50820 81564
rect 81276 81508 81332 81564
rect 81380 81508 81436 81564
rect 81484 81508 81540 81564
rect 4476 80724 4532 80780
rect 4580 80724 4636 80780
rect 4684 80724 4740 80780
rect 35196 80724 35252 80780
rect 35300 80724 35356 80780
rect 35404 80724 35460 80780
rect 65916 80724 65972 80780
rect 66020 80724 66076 80780
rect 66124 80724 66180 80780
rect 96636 80724 96692 80780
rect 96740 80724 96796 80780
rect 96844 80724 96900 80780
rect 19836 79940 19892 79996
rect 19940 79940 19996 79996
rect 20044 79940 20100 79996
rect 50556 79940 50612 79996
rect 50660 79940 50716 79996
rect 50764 79940 50820 79996
rect 81276 79940 81332 79996
rect 81380 79940 81436 79996
rect 81484 79940 81540 79996
rect 4476 79156 4532 79212
rect 4580 79156 4636 79212
rect 4684 79156 4740 79212
rect 35196 79156 35252 79212
rect 35300 79156 35356 79212
rect 35404 79156 35460 79212
rect 65916 79156 65972 79212
rect 66020 79156 66076 79212
rect 66124 79156 66180 79212
rect 96636 79156 96692 79212
rect 96740 79156 96796 79212
rect 96844 79156 96900 79212
rect 19836 78372 19892 78428
rect 19940 78372 19996 78428
rect 20044 78372 20100 78428
rect 50556 78372 50612 78428
rect 50660 78372 50716 78428
rect 50764 78372 50820 78428
rect 81276 78372 81332 78428
rect 81380 78372 81436 78428
rect 81484 78372 81540 78428
rect 4476 77588 4532 77644
rect 4580 77588 4636 77644
rect 4684 77588 4740 77644
rect 35196 77588 35252 77644
rect 35300 77588 35356 77644
rect 35404 77588 35460 77644
rect 65916 77588 65972 77644
rect 66020 77588 66076 77644
rect 66124 77588 66180 77644
rect 96636 77588 96692 77644
rect 96740 77588 96796 77644
rect 96844 77588 96900 77644
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 81276 76804 81332 76860
rect 81380 76804 81436 76860
rect 81484 76804 81540 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 96636 76020 96692 76076
rect 96740 76020 96796 76076
rect 96844 76020 96900 76076
rect 71932 75740 71988 75796
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 81276 75236 81332 75292
rect 81380 75236 81436 75292
rect 81484 75236 81540 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 96636 74452 96692 74508
rect 96740 74452 96796 74508
rect 96844 74452 96900 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 81276 73668 81332 73724
rect 81380 73668 81436 73724
rect 81484 73668 81540 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 96636 72884 96692 72940
rect 96740 72884 96796 72940
rect 96844 72884 96900 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 81276 72100 81332 72156
rect 81380 72100 81436 72156
rect 81484 72100 81540 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 96636 71316 96692 71372
rect 96740 71316 96796 71372
rect 96844 71316 96900 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 81276 70532 81332 70588
rect 81380 70532 81436 70588
rect 81484 70532 81540 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 96636 69748 96692 69804
rect 96740 69748 96796 69804
rect 96844 69748 96900 69804
rect 76300 69468 76356 69524
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 81276 68964 81332 69020
rect 81380 68964 81436 69020
rect 81484 68964 81540 69020
rect 73388 68684 73444 68740
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 96636 68180 96692 68236
rect 96740 68180 96796 68236
rect 96844 68180 96900 68236
rect 71372 68124 71428 68180
rect 76300 67676 76356 67732
rect 71596 67564 71652 67620
rect 74508 67452 74564 67508
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 81276 67396 81332 67452
rect 81380 67396 81436 67452
rect 81484 67396 81540 67452
rect 73388 67340 73444 67396
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 96636 66612 96692 66668
rect 96740 66612 96796 66668
rect 96844 66612 96900 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 81276 65828 81332 65884
rect 81380 65828 81436 65884
rect 81484 65828 81540 65884
rect 82796 65100 82852 65156
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 96636 65044 96692 65100
rect 96740 65044 96796 65100
rect 96844 65044 96900 65100
rect 82908 64988 82964 65044
rect 70700 64876 70756 64932
rect 71596 64652 71652 64708
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 81276 64260 81332 64316
rect 81380 64260 81436 64316
rect 81484 64260 81540 64316
rect 79660 64204 79716 64260
rect 72940 64092 72996 64148
rect 70700 63980 70756 64036
rect 82796 63980 82852 64036
rect 72940 63868 72996 63924
rect 82908 63756 82964 63812
rect 82796 63644 82852 63700
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 96636 63476 96692 63532
rect 96740 63476 96796 63532
rect 96844 63476 96900 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 81276 62692 81332 62748
rect 81380 62692 81436 62748
rect 81484 62692 81540 62748
rect 83580 62412 83636 62468
rect 74508 62300 74564 62356
rect 83692 62300 83748 62356
rect 71372 62188 71428 62244
rect 83580 62076 83636 62132
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 96636 61908 96692 61964
rect 96740 61908 96796 61964
rect 96844 61908 96900 61964
rect 83580 61516 83636 61572
rect 79660 61292 79716 61348
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 81276 61124 81332 61180
rect 81380 61124 81436 61180
rect 81484 61124 81540 61180
rect 85596 60620 85652 60676
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 96636 60340 96692 60396
rect 96740 60340 96796 60396
rect 96844 60340 96900 60396
rect 79660 60284 79716 60340
rect 71932 60172 71988 60228
rect 71932 59948 71988 60004
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 81276 59556 81332 59612
rect 81380 59556 81436 59612
rect 81484 59556 81540 59612
rect 83692 59500 83748 59556
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 96636 58772 96692 58828
rect 96740 58772 96796 58828
rect 96844 58772 96900 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 81276 57988 81332 58044
rect 81380 57988 81436 58044
rect 81484 57988 81540 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 96636 57204 96692 57260
rect 96740 57204 96796 57260
rect 96844 57204 96900 57260
rect 74956 57148 75012 57204
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 81276 56420 81332 56476
rect 81380 56420 81436 56476
rect 81484 56420 81540 56476
rect 85596 56252 85652 56308
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 96636 55636 96692 55692
rect 96740 55636 96796 55692
rect 96844 55636 96900 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 81276 54852 81332 54908
rect 81380 54852 81436 54908
rect 81484 54852 81540 54908
rect 90860 54572 90916 54628
rect 90860 54348 90916 54404
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 96636 54068 96692 54124
rect 96740 54068 96796 54124
rect 96844 54068 96900 54124
rect 93660 54012 93716 54068
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 81276 53284 81332 53340
rect 81380 53284 81436 53340
rect 81484 53284 81540 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 96636 52500 96692 52556
rect 96740 52500 96796 52556
rect 96844 52500 96900 52556
rect 93660 51772 93716 51828
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 81276 51716 81332 51772
rect 81380 51716 81436 51772
rect 81484 51716 81540 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 96636 50932 96692 50988
rect 96740 50932 96796 50988
rect 96844 50932 96900 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 81276 50148 81332 50204
rect 81380 50148 81436 50204
rect 81484 50148 81540 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 96636 49364 96692 49420
rect 96740 49364 96796 49420
rect 96844 49364 96900 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 81276 48580 81332 48636
rect 81380 48580 81436 48636
rect 81484 48580 81540 48636
rect 74956 48524 75012 48580
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 96636 47796 96692 47852
rect 96740 47796 96796 47852
rect 96844 47796 96900 47852
rect 94220 47404 94276 47460
rect 94220 47068 94276 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 81276 47012 81332 47068
rect 81380 47012 81436 47068
rect 81484 47012 81540 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
<< metal4 >>
rect 4448 96460 4768 96492
rect 4448 96404 4476 96460
rect 4532 96404 4580 96460
rect 4636 96404 4684 96460
rect 4740 96404 4768 96460
rect 4448 94892 4768 96404
rect 4448 94836 4476 94892
rect 4532 94836 4580 94892
rect 4636 94836 4684 94892
rect 4740 94836 4768 94892
rect 4448 93324 4768 94836
rect 4448 93268 4476 93324
rect 4532 93268 4580 93324
rect 4636 93268 4684 93324
rect 4740 93268 4768 93324
rect 4448 91756 4768 93268
rect 4448 91700 4476 91756
rect 4532 91700 4580 91756
rect 4636 91700 4684 91756
rect 4740 91700 4768 91756
rect 4448 90188 4768 91700
rect 4448 90132 4476 90188
rect 4532 90132 4580 90188
rect 4636 90132 4684 90188
rect 4740 90132 4768 90188
rect 4448 88620 4768 90132
rect 4448 88564 4476 88620
rect 4532 88564 4580 88620
rect 4636 88564 4684 88620
rect 4740 88564 4768 88620
rect 4448 87052 4768 88564
rect 4448 86996 4476 87052
rect 4532 86996 4580 87052
rect 4636 86996 4684 87052
rect 4740 86996 4768 87052
rect 4448 85484 4768 86996
rect 4448 85428 4476 85484
rect 4532 85428 4580 85484
rect 4636 85428 4684 85484
rect 4740 85428 4768 85484
rect 4448 83916 4768 85428
rect 4448 83860 4476 83916
rect 4532 83860 4580 83916
rect 4636 83860 4684 83916
rect 4740 83860 4768 83916
rect 4448 82348 4768 83860
rect 4448 82292 4476 82348
rect 4532 82292 4580 82348
rect 4636 82292 4684 82348
rect 4740 82292 4768 82348
rect 4448 80780 4768 82292
rect 4448 80724 4476 80780
rect 4532 80724 4580 80780
rect 4636 80724 4684 80780
rect 4740 80724 4768 80780
rect 4448 79212 4768 80724
rect 4448 79156 4476 79212
rect 4532 79156 4580 79212
rect 4636 79156 4684 79212
rect 4740 79156 4768 79212
rect 4448 77644 4768 79156
rect 4448 77588 4476 77644
rect 4532 77588 4580 77644
rect 4636 77588 4684 77644
rect 4740 77588 4768 77644
rect 4448 76076 4768 77588
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 95676 20128 96492
rect 19808 95620 19836 95676
rect 19892 95620 19940 95676
rect 19996 95620 20044 95676
rect 20100 95620 20128 95676
rect 19808 94108 20128 95620
rect 19808 94052 19836 94108
rect 19892 94052 19940 94108
rect 19996 94052 20044 94108
rect 20100 94052 20128 94108
rect 19808 92540 20128 94052
rect 19808 92484 19836 92540
rect 19892 92484 19940 92540
rect 19996 92484 20044 92540
rect 20100 92484 20128 92540
rect 19808 90972 20128 92484
rect 19808 90916 19836 90972
rect 19892 90916 19940 90972
rect 19996 90916 20044 90972
rect 20100 90916 20128 90972
rect 19808 89404 20128 90916
rect 19808 89348 19836 89404
rect 19892 89348 19940 89404
rect 19996 89348 20044 89404
rect 20100 89348 20128 89404
rect 19808 87836 20128 89348
rect 19808 87780 19836 87836
rect 19892 87780 19940 87836
rect 19996 87780 20044 87836
rect 20100 87780 20128 87836
rect 19808 86268 20128 87780
rect 19808 86212 19836 86268
rect 19892 86212 19940 86268
rect 19996 86212 20044 86268
rect 20100 86212 20128 86268
rect 19808 84700 20128 86212
rect 19808 84644 19836 84700
rect 19892 84644 19940 84700
rect 19996 84644 20044 84700
rect 20100 84644 20128 84700
rect 19808 83132 20128 84644
rect 19808 83076 19836 83132
rect 19892 83076 19940 83132
rect 19996 83076 20044 83132
rect 20100 83076 20128 83132
rect 19808 81564 20128 83076
rect 19808 81508 19836 81564
rect 19892 81508 19940 81564
rect 19996 81508 20044 81564
rect 20100 81508 20128 81564
rect 19808 79996 20128 81508
rect 19808 79940 19836 79996
rect 19892 79940 19940 79996
rect 19996 79940 20044 79996
rect 20100 79940 20128 79996
rect 19808 78428 20128 79940
rect 19808 78372 19836 78428
rect 19892 78372 19940 78428
rect 19996 78372 20044 78428
rect 20100 78372 20128 78428
rect 19808 76860 20128 78372
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 96460 35488 96492
rect 35168 96404 35196 96460
rect 35252 96404 35300 96460
rect 35356 96404 35404 96460
rect 35460 96404 35488 96460
rect 35168 94892 35488 96404
rect 35168 94836 35196 94892
rect 35252 94836 35300 94892
rect 35356 94836 35404 94892
rect 35460 94836 35488 94892
rect 35168 93324 35488 94836
rect 35168 93268 35196 93324
rect 35252 93268 35300 93324
rect 35356 93268 35404 93324
rect 35460 93268 35488 93324
rect 35168 91756 35488 93268
rect 35168 91700 35196 91756
rect 35252 91700 35300 91756
rect 35356 91700 35404 91756
rect 35460 91700 35488 91756
rect 35168 90188 35488 91700
rect 35168 90132 35196 90188
rect 35252 90132 35300 90188
rect 35356 90132 35404 90188
rect 35460 90132 35488 90188
rect 35168 88620 35488 90132
rect 35168 88564 35196 88620
rect 35252 88564 35300 88620
rect 35356 88564 35404 88620
rect 35460 88564 35488 88620
rect 35168 87052 35488 88564
rect 35168 86996 35196 87052
rect 35252 86996 35300 87052
rect 35356 86996 35404 87052
rect 35460 86996 35488 87052
rect 35168 85484 35488 86996
rect 35168 85428 35196 85484
rect 35252 85428 35300 85484
rect 35356 85428 35404 85484
rect 35460 85428 35488 85484
rect 35168 83916 35488 85428
rect 35168 83860 35196 83916
rect 35252 83860 35300 83916
rect 35356 83860 35404 83916
rect 35460 83860 35488 83916
rect 35168 82348 35488 83860
rect 35168 82292 35196 82348
rect 35252 82292 35300 82348
rect 35356 82292 35404 82348
rect 35460 82292 35488 82348
rect 35168 80780 35488 82292
rect 35168 80724 35196 80780
rect 35252 80724 35300 80780
rect 35356 80724 35404 80780
rect 35460 80724 35488 80780
rect 35168 79212 35488 80724
rect 35168 79156 35196 79212
rect 35252 79156 35300 79212
rect 35356 79156 35404 79212
rect 35460 79156 35488 79212
rect 35168 77644 35488 79156
rect 35168 77588 35196 77644
rect 35252 77588 35300 77644
rect 35356 77588 35404 77644
rect 35460 77588 35488 77644
rect 35168 76076 35488 77588
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 95676 50848 96492
rect 50528 95620 50556 95676
rect 50612 95620 50660 95676
rect 50716 95620 50764 95676
rect 50820 95620 50848 95676
rect 50528 94108 50848 95620
rect 50528 94052 50556 94108
rect 50612 94052 50660 94108
rect 50716 94052 50764 94108
rect 50820 94052 50848 94108
rect 50528 92540 50848 94052
rect 50528 92484 50556 92540
rect 50612 92484 50660 92540
rect 50716 92484 50764 92540
rect 50820 92484 50848 92540
rect 50528 90972 50848 92484
rect 50528 90916 50556 90972
rect 50612 90916 50660 90972
rect 50716 90916 50764 90972
rect 50820 90916 50848 90972
rect 50528 89404 50848 90916
rect 50528 89348 50556 89404
rect 50612 89348 50660 89404
rect 50716 89348 50764 89404
rect 50820 89348 50848 89404
rect 50528 87836 50848 89348
rect 50528 87780 50556 87836
rect 50612 87780 50660 87836
rect 50716 87780 50764 87836
rect 50820 87780 50848 87836
rect 50528 86268 50848 87780
rect 50528 86212 50556 86268
rect 50612 86212 50660 86268
rect 50716 86212 50764 86268
rect 50820 86212 50848 86268
rect 50528 84700 50848 86212
rect 50528 84644 50556 84700
rect 50612 84644 50660 84700
rect 50716 84644 50764 84700
rect 50820 84644 50848 84700
rect 50528 83132 50848 84644
rect 50528 83076 50556 83132
rect 50612 83076 50660 83132
rect 50716 83076 50764 83132
rect 50820 83076 50848 83132
rect 50528 81564 50848 83076
rect 50528 81508 50556 81564
rect 50612 81508 50660 81564
rect 50716 81508 50764 81564
rect 50820 81508 50848 81564
rect 50528 79996 50848 81508
rect 50528 79940 50556 79996
rect 50612 79940 50660 79996
rect 50716 79940 50764 79996
rect 50820 79940 50848 79996
rect 50528 78428 50848 79940
rect 50528 78372 50556 78428
rect 50612 78372 50660 78428
rect 50716 78372 50764 78428
rect 50820 78372 50848 78428
rect 50528 76860 50848 78372
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 96460 66208 96492
rect 65888 96404 65916 96460
rect 65972 96404 66020 96460
rect 66076 96404 66124 96460
rect 66180 96404 66208 96460
rect 65888 94892 66208 96404
rect 65888 94836 65916 94892
rect 65972 94836 66020 94892
rect 66076 94836 66124 94892
rect 66180 94836 66208 94892
rect 65888 93324 66208 94836
rect 65888 93268 65916 93324
rect 65972 93268 66020 93324
rect 66076 93268 66124 93324
rect 66180 93268 66208 93324
rect 65888 91756 66208 93268
rect 65888 91700 65916 91756
rect 65972 91700 66020 91756
rect 66076 91700 66124 91756
rect 66180 91700 66208 91756
rect 65888 90188 66208 91700
rect 65888 90132 65916 90188
rect 65972 90132 66020 90188
rect 66076 90132 66124 90188
rect 66180 90132 66208 90188
rect 65888 88620 66208 90132
rect 65888 88564 65916 88620
rect 65972 88564 66020 88620
rect 66076 88564 66124 88620
rect 66180 88564 66208 88620
rect 65888 87052 66208 88564
rect 65888 86996 65916 87052
rect 65972 86996 66020 87052
rect 66076 86996 66124 87052
rect 66180 86996 66208 87052
rect 65888 85484 66208 86996
rect 65888 85428 65916 85484
rect 65972 85428 66020 85484
rect 66076 85428 66124 85484
rect 66180 85428 66208 85484
rect 65888 83916 66208 85428
rect 65888 83860 65916 83916
rect 65972 83860 66020 83916
rect 66076 83860 66124 83916
rect 66180 83860 66208 83916
rect 65888 82348 66208 83860
rect 65888 82292 65916 82348
rect 65972 82292 66020 82348
rect 66076 82292 66124 82348
rect 66180 82292 66208 82348
rect 65888 80780 66208 82292
rect 65888 80724 65916 80780
rect 65972 80724 66020 80780
rect 66076 80724 66124 80780
rect 66180 80724 66208 80780
rect 65888 79212 66208 80724
rect 65888 79156 65916 79212
rect 65972 79156 66020 79212
rect 66076 79156 66124 79212
rect 66180 79156 66208 79212
rect 65888 77644 66208 79156
rect 65888 77588 65916 77644
rect 65972 77588 66020 77644
rect 66076 77588 66124 77644
rect 66180 77588 66208 77644
rect 65888 76076 66208 77588
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 81248 95676 81568 96492
rect 81248 95620 81276 95676
rect 81332 95620 81380 95676
rect 81436 95620 81484 95676
rect 81540 95620 81568 95676
rect 81248 94108 81568 95620
rect 81248 94052 81276 94108
rect 81332 94052 81380 94108
rect 81436 94052 81484 94108
rect 81540 94052 81568 94108
rect 81248 92540 81568 94052
rect 81248 92484 81276 92540
rect 81332 92484 81380 92540
rect 81436 92484 81484 92540
rect 81540 92484 81568 92540
rect 81248 90972 81568 92484
rect 81248 90916 81276 90972
rect 81332 90916 81380 90972
rect 81436 90916 81484 90972
rect 81540 90916 81568 90972
rect 81248 89404 81568 90916
rect 81248 89348 81276 89404
rect 81332 89348 81380 89404
rect 81436 89348 81484 89404
rect 81540 89348 81568 89404
rect 81248 87836 81568 89348
rect 81248 87780 81276 87836
rect 81332 87780 81380 87836
rect 81436 87780 81484 87836
rect 81540 87780 81568 87836
rect 81248 86268 81568 87780
rect 81248 86212 81276 86268
rect 81332 86212 81380 86268
rect 81436 86212 81484 86268
rect 81540 86212 81568 86268
rect 81248 84700 81568 86212
rect 81248 84644 81276 84700
rect 81332 84644 81380 84700
rect 81436 84644 81484 84700
rect 81540 84644 81568 84700
rect 81248 83132 81568 84644
rect 81248 83076 81276 83132
rect 81332 83076 81380 83132
rect 81436 83076 81484 83132
rect 81540 83076 81568 83132
rect 81248 81564 81568 83076
rect 81248 81508 81276 81564
rect 81332 81508 81380 81564
rect 81436 81508 81484 81564
rect 81540 81508 81568 81564
rect 81248 79996 81568 81508
rect 81248 79940 81276 79996
rect 81332 79940 81380 79996
rect 81436 79940 81484 79996
rect 81540 79940 81568 79996
rect 81248 78428 81568 79940
rect 81248 78372 81276 78428
rect 81332 78372 81380 78428
rect 81436 78372 81484 78428
rect 81540 78372 81568 78428
rect 81248 76860 81568 78372
rect 81248 76804 81276 76860
rect 81332 76804 81380 76860
rect 81436 76804 81484 76860
rect 81540 76804 81568 76860
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 71932 75796 71988 75806
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 71372 68180 71428 68190
rect 70700 64932 70756 64942
rect 70700 64036 70756 64876
rect 70700 63970 70756 63980
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 71372 62244 71428 68124
rect 71596 67620 71652 67630
rect 71596 64708 71652 67564
rect 71596 64642 71652 64652
rect 71372 62178 71428 62188
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 71932 60228 71988 75740
rect 81248 75292 81568 76804
rect 81248 75236 81276 75292
rect 81332 75236 81380 75292
rect 81436 75236 81484 75292
rect 81540 75236 81568 75292
rect 81248 73724 81568 75236
rect 81248 73668 81276 73724
rect 81332 73668 81380 73724
rect 81436 73668 81484 73724
rect 81540 73668 81568 73724
rect 81248 72156 81568 73668
rect 81248 72100 81276 72156
rect 81332 72100 81380 72156
rect 81436 72100 81484 72156
rect 81540 72100 81568 72156
rect 81248 70588 81568 72100
rect 81248 70532 81276 70588
rect 81332 70532 81380 70588
rect 81436 70532 81484 70588
rect 81540 70532 81568 70588
rect 76300 69524 76356 69534
rect 73388 68740 73444 68750
rect 73388 67396 73444 68684
rect 76300 67732 76356 69468
rect 76300 67666 76356 67676
rect 81248 69020 81568 70532
rect 81248 68964 81276 69020
rect 81332 68964 81380 69020
rect 81436 68964 81484 69020
rect 81540 68964 81568 69020
rect 73388 67330 73444 67340
rect 74508 67508 74564 67518
rect 72940 64148 72996 64158
rect 72940 63924 72996 64092
rect 72940 63858 72996 63868
rect 74508 62356 74564 67452
rect 81248 67452 81568 68964
rect 81248 67396 81276 67452
rect 81332 67396 81380 67452
rect 81436 67396 81484 67452
rect 81540 67396 81568 67452
rect 81248 65884 81568 67396
rect 81248 65828 81276 65884
rect 81332 65828 81380 65884
rect 81436 65828 81484 65884
rect 81540 65828 81568 65884
rect 81248 64316 81568 65828
rect 96608 96460 96928 96492
rect 96608 96404 96636 96460
rect 96692 96404 96740 96460
rect 96796 96404 96844 96460
rect 96900 96404 96928 96460
rect 96608 94892 96928 96404
rect 96608 94836 96636 94892
rect 96692 94836 96740 94892
rect 96796 94836 96844 94892
rect 96900 94836 96928 94892
rect 96608 93324 96928 94836
rect 96608 93268 96636 93324
rect 96692 93268 96740 93324
rect 96796 93268 96844 93324
rect 96900 93268 96928 93324
rect 96608 91756 96928 93268
rect 96608 91700 96636 91756
rect 96692 91700 96740 91756
rect 96796 91700 96844 91756
rect 96900 91700 96928 91756
rect 96608 90188 96928 91700
rect 96608 90132 96636 90188
rect 96692 90132 96740 90188
rect 96796 90132 96844 90188
rect 96900 90132 96928 90188
rect 96608 88620 96928 90132
rect 96608 88564 96636 88620
rect 96692 88564 96740 88620
rect 96796 88564 96844 88620
rect 96900 88564 96928 88620
rect 96608 87052 96928 88564
rect 96608 86996 96636 87052
rect 96692 86996 96740 87052
rect 96796 86996 96844 87052
rect 96900 86996 96928 87052
rect 96608 85484 96928 86996
rect 96608 85428 96636 85484
rect 96692 85428 96740 85484
rect 96796 85428 96844 85484
rect 96900 85428 96928 85484
rect 96608 83916 96928 85428
rect 96608 83860 96636 83916
rect 96692 83860 96740 83916
rect 96796 83860 96844 83916
rect 96900 83860 96928 83916
rect 96608 82348 96928 83860
rect 96608 82292 96636 82348
rect 96692 82292 96740 82348
rect 96796 82292 96844 82348
rect 96900 82292 96928 82348
rect 96608 80780 96928 82292
rect 96608 80724 96636 80780
rect 96692 80724 96740 80780
rect 96796 80724 96844 80780
rect 96900 80724 96928 80780
rect 96608 79212 96928 80724
rect 96608 79156 96636 79212
rect 96692 79156 96740 79212
rect 96796 79156 96844 79212
rect 96900 79156 96928 79212
rect 96608 77644 96928 79156
rect 96608 77588 96636 77644
rect 96692 77588 96740 77644
rect 96796 77588 96844 77644
rect 96900 77588 96928 77644
rect 96608 76076 96928 77588
rect 96608 76020 96636 76076
rect 96692 76020 96740 76076
rect 96796 76020 96844 76076
rect 96900 76020 96928 76076
rect 96608 74508 96928 76020
rect 96608 74452 96636 74508
rect 96692 74452 96740 74508
rect 96796 74452 96844 74508
rect 96900 74452 96928 74508
rect 96608 72940 96928 74452
rect 96608 72884 96636 72940
rect 96692 72884 96740 72940
rect 96796 72884 96844 72940
rect 96900 72884 96928 72940
rect 96608 71372 96928 72884
rect 96608 71316 96636 71372
rect 96692 71316 96740 71372
rect 96796 71316 96844 71372
rect 96900 71316 96928 71372
rect 96608 69804 96928 71316
rect 96608 69748 96636 69804
rect 96692 69748 96740 69804
rect 96796 69748 96844 69804
rect 96900 69748 96928 69804
rect 96608 68236 96928 69748
rect 96608 68180 96636 68236
rect 96692 68180 96740 68236
rect 96796 68180 96844 68236
rect 96900 68180 96928 68236
rect 96608 66668 96928 68180
rect 96608 66612 96636 66668
rect 96692 66612 96740 66668
rect 96796 66612 96844 66668
rect 96900 66612 96928 66668
rect 74508 62290 74564 62300
rect 79660 64260 79716 64270
rect 79660 61348 79716 64204
rect 79660 60340 79716 61292
rect 79660 60274 79716 60284
rect 81248 64260 81276 64316
rect 81332 64260 81380 64316
rect 81436 64260 81484 64316
rect 81540 64260 81568 64316
rect 81248 62748 81568 64260
rect 82796 65156 82852 65166
rect 82796 64036 82852 65100
rect 96608 65100 96928 66612
rect 82796 63700 82852 63980
rect 82908 65044 82964 65054
rect 82908 63812 82964 64988
rect 82908 63746 82964 63756
rect 96608 65044 96636 65100
rect 96692 65044 96740 65100
rect 96796 65044 96844 65100
rect 96900 65044 96928 65100
rect 82796 63634 82852 63644
rect 81248 62692 81276 62748
rect 81332 62692 81380 62748
rect 81436 62692 81484 62748
rect 81540 62692 81568 62748
rect 81248 61180 81568 62692
rect 96608 63532 96928 65044
rect 96608 63476 96636 63532
rect 96692 63476 96740 63532
rect 96796 63476 96844 63532
rect 96900 63476 96928 63532
rect 83580 62468 83636 62478
rect 83580 62132 83636 62412
rect 83580 61572 83636 62076
rect 83580 61506 83636 61516
rect 83692 62356 83748 62366
rect 81248 61124 81276 61180
rect 81332 61124 81380 61180
rect 81436 61124 81484 61180
rect 81540 61124 81568 61180
rect 71932 60004 71988 60172
rect 71932 59938 71988 59948
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 81248 59612 81568 61124
rect 81248 59556 81276 59612
rect 81332 59556 81380 59612
rect 81436 59556 81484 59612
rect 81540 59556 81568 59612
rect 81248 58044 81568 59556
rect 83692 59556 83748 62300
rect 96608 61964 96928 63476
rect 96608 61908 96636 61964
rect 96692 61908 96740 61964
rect 96796 61908 96844 61964
rect 96900 61908 96928 61964
rect 83692 59490 83748 59500
rect 85596 60676 85652 60686
rect 81248 57988 81276 58044
rect 81332 57988 81380 58044
rect 81436 57988 81484 58044
rect 81540 57988 81568 58044
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 74956 57204 75012 57214
rect 74956 48580 75012 57148
rect 74956 48514 75012 48524
rect 81248 56476 81568 57988
rect 81248 56420 81276 56476
rect 81332 56420 81380 56476
rect 81436 56420 81484 56476
rect 81540 56420 81568 56476
rect 81248 54908 81568 56420
rect 85596 56308 85652 60620
rect 85596 56242 85652 56252
rect 96608 60396 96928 61908
rect 96608 60340 96636 60396
rect 96692 60340 96740 60396
rect 96796 60340 96844 60396
rect 96900 60340 96928 60396
rect 96608 58828 96928 60340
rect 96608 58772 96636 58828
rect 96692 58772 96740 58828
rect 96796 58772 96844 58828
rect 96900 58772 96928 58828
rect 96608 57260 96928 58772
rect 96608 57204 96636 57260
rect 96692 57204 96740 57260
rect 96796 57204 96844 57260
rect 96900 57204 96928 57260
rect 81248 54852 81276 54908
rect 81332 54852 81380 54908
rect 81436 54852 81484 54908
rect 81540 54852 81568 54908
rect 81248 53340 81568 54852
rect 96608 55692 96928 57204
rect 96608 55636 96636 55692
rect 96692 55636 96740 55692
rect 96796 55636 96844 55692
rect 96900 55636 96928 55692
rect 90860 54628 90916 54638
rect 90860 54404 90916 54572
rect 90860 54338 90916 54348
rect 96608 54124 96928 55636
rect 81248 53284 81276 53340
rect 81332 53284 81380 53340
rect 81436 53284 81484 53340
rect 81540 53284 81568 53340
rect 81248 51772 81568 53284
rect 81248 51716 81276 51772
rect 81332 51716 81380 51772
rect 81436 51716 81484 51772
rect 81540 51716 81568 51772
rect 93660 54068 93716 54078
rect 93660 51828 93716 54012
rect 93660 51762 93716 51772
rect 96608 54068 96636 54124
rect 96692 54068 96740 54124
rect 96796 54068 96844 54124
rect 96900 54068 96928 54124
rect 96608 52556 96928 54068
rect 96608 52500 96636 52556
rect 96692 52500 96740 52556
rect 96796 52500 96844 52556
rect 96900 52500 96928 52556
rect 81248 50204 81568 51716
rect 81248 50148 81276 50204
rect 81332 50148 81380 50204
rect 81436 50148 81484 50204
rect 81540 50148 81568 50204
rect 81248 48636 81568 50148
rect 81248 48580 81276 48636
rect 81332 48580 81380 48636
rect 81436 48580 81484 48636
rect 81540 48580 81568 48636
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 81248 47068 81568 48580
rect 96608 50988 96928 52500
rect 96608 50932 96636 50988
rect 96692 50932 96740 50988
rect 96796 50932 96844 50988
rect 96900 50932 96928 50988
rect 96608 49420 96928 50932
rect 96608 49364 96636 49420
rect 96692 49364 96740 49420
rect 96796 49364 96844 49420
rect 96900 49364 96928 49420
rect 96608 47852 96928 49364
rect 96608 47796 96636 47852
rect 96692 47796 96740 47852
rect 96796 47796 96844 47852
rect 96900 47796 96928 47852
rect 81248 47012 81276 47068
rect 81332 47012 81380 47068
rect 81436 47012 81484 47068
rect 81540 47012 81568 47068
rect 94220 47460 94276 47470
rect 94220 47124 94276 47404
rect 94220 47058 94276 47068
rect 81248 45500 81568 47012
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 81248 21980 81568 23492
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 81248 17276 81568 18788
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 81248 15708 81568 17220
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 81248 12572 81568 14084
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 81248 11004 81568 12516
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 81248 7868 81568 9380
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 81248 6300 81568 7812
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 81248 4732 81568 6244
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 81248 3164 81568 4676
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 96608 46284 96928 47796
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 96608 19628 96928 21140
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0831__I pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 70560 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__I
timestamp 1669390400
transform 1 0 81872 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__I
timestamp 1669390400
transform 1 0 68432 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__I
timestamp 1669390400
transform 1 0 78512 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__I0
timestamp 1669390400
transform -1 0 80304 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__S0
timestamp 1669390400
transform 1 0 80752 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__S1
timestamp 1669390400
transform -1 0 80528 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__A1
timestamp 1669390400
transform 1 0 82768 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__A2
timestamp 1669390400
transform 1 0 82320 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0841__I
timestamp 1669390400
transform 1 0 72576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__I
timestamp 1669390400
transform 1 0 82768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__I
timestamp 1669390400
transform -1 0 82768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0845__I
timestamp 1669390400
transform 1 0 66192 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0846__I
timestamp 1669390400
transform 1 0 82992 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__I1
timestamp 1669390400
transform 1 0 84336 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__I2
timestamp 1669390400
transform 1 0 82320 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__S0
timestamp 1669390400
transform -1 0 82992 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__S1
timestamp 1669390400
transform -1 0 81872 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__I
timestamp 1669390400
transform 1 0 69216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__I
timestamp 1669390400
transform 1 0 71232 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__I
timestamp 1669390400
transform 1 0 83216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__B
timestamp 1669390400
transform 1 0 85120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__I
timestamp 1669390400
transform -1 0 82320 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0853__I
timestamp 1669390400
transform 1 0 73024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__I
timestamp 1669390400
transform 1 0 75712 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0856__I
timestamp 1669390400
transform 1 0 77392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__I2
timestamp 1669390400
transform 1 0 76944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__S0
timestamp 1669390400
transform -1 0 77616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__S1
timestamp 1669390400
transform -1 0 78288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A1
timestamp 1669390400
transform 1 0 83552 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A2
timestamp 1669390400
transform 1 0 84336 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__I
timestamp 1669390400
transform 1 0 70336 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__I
timestamp 1669390400
transform 1 0 71232 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__I
timestamp 1669390400
transform 1 0 82544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__I0
timestamp 1669390400
transform 1 0 83888 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__I1
timestamp 1669390400
transform 1 0 84336 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__I3
timestamp 1669390400
transform 1 0 84448 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__S0
timestamp 1669390400
transform 1 0 83104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__S1
timestamp 1669390400
transform 1 0 83440 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__I
timestamp 1669390400
transform 1 0 71344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__I
timestamp 1669390400
transform 1 0 81200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A1
timestamp 1669390400
transform -1 0 83216 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__I0
timestamp 1669390400
transform -1 0 89600 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__S0
timestamp 1669390400
transform 1 0 86464 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0869__S1
timestamp 1669390400
transform 1 0 86016 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A1
timestamp 1669390400
transform 1 0 87024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A2
timestamp 1669390400
transform 1 0 86464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__I1
timestamp 1669390400
transform -1 0 93296 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__I2
timestamp 1669390400
transform -1 0 93184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__S0
timestamp 1669390400
transform 1 0 89152 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__S1
timestamp 1669390400
transform -1 0 88928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__B
timestamp 1669390400
transform 1 0 87920 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__I1
timestamp 1669390400
transform -1 0 88704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__I2
timestamp 1669390400
transform 1 0 89040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__S0
timestamp 1669390400
transform -1 0 85232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__S1
timestamp 1669390400
transform -1 0 84224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__A1
timestamp 1669390400
transform -1 0 84224 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__A2
timestamp 1669390400
transform 1 0 85680 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__I0
timestamp 1669390400
transform -1 0 89376 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__I1
timestamp 1669390400
transform -1 0 89824 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__I3
timestamp 1669390400
transform 1 0 88480 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__S0
timestamp 1669390400
transform 1 0 85120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__S1
timestamp 1669390400
transform 1 0 84448 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__A1
timestamp 1669390400
transform 1 0 86912 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__I
timestamp 1669390400
transform 1 0 71008 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__I0
timestamp 1669390400
transform 1 0 89600 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__S0
timestamp 1669390400
transform -1 0 85904 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__S1
timestamp 1669390400
transform 1 0 89152 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__A1
timestamp 1669390400
transform 1 0 83552 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__A2
timestamp 1669390400
transform 1 0 85120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__I1
timestamp 1669390400
transform 1 0 93408 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__I2
timestamp 1669390400
transform 1 0 92960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__S0
timestamp 1669390400
transform 1 0 89600 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__S1
timestamp 1669390400
transform 1 0 91168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0884__B
timestamp 1669390400
transform -1 0 87472 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__I0
timestamp 1669390400
transform 1 0 90384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__I3
timestamp 1669390400
transform -1 0 89712 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__S0
timestamp 1669390400
transform 1 0 85680 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__S1
timestamp 1669390400
transform 1 0 85456 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A1
timestamp 1669390400
transform 1 0 87024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0886__A2
timestamp 1669390400
transform 1 0 87472 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__I
timestamp 1669390400
transform 1 0 85120 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__I
timestamp 1669390400
transform -1 0 69664 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I1
timestamp 1669390400
transform -1 0 87584 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I2
timestamp 1669390400
transform 1 0 87360 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I3
timestamp 1669390400
transform -1 0 87360 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__S0
timestamp 1669390400
transform 1 0 83104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__S1
timestamp 1669390400
transform 1 0 83552 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0890__A1
timestamp 1669390400
transform 1 0 86240 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__S0
timestamp 1669390400
transform 1 0 86128 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__S1
timestamp 1669390400
transform -1 0 85792 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A1
timestamp 1669390400
transform 1 0 88256 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A2
timestamp 1669390400
transform 1 0 87024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__I1
timestamp 1669390400
transform 1 0 92176 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__I2
timestamp 1669390400
transform 1 0 91728 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__S0
timestamp 1669390400
transform 1 0 88256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__S1
timestamp 1669390400
transform 1 0 88368 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0895__B
timestamp 1669390400
transform 1 0 87360 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__I0
timestamp 1669390400
transform 1 0 85008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__I1
timestamp 1669390400
transform 1 0 85456 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__I2
timestamp 1669390400
transform 1 0 85232 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__S0
timestamp 1669390400
transform 1 0 80976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__S1
timestamp 1669390400
transform 1 0 80528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A1
timestamp 1669390400
transform 1 0 87136 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A2
timestamp 1669390400
transform 1 0 86688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__I0
timestamp 1669390400
transform 1 0 89376 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__I1
timestamp 1669390400
transform 1 0 89824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__I3
timestamp 1669390400
transform -1 0 89152 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__S0
timestamp 1669390400
transform 1 0 84784 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__S1
timestamp 1669390400
transform 1 0 85232 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__A1
timestamp 1669390400
transform 1 0 87584 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__I
timestamp 1669390400
transform 1 0 68432 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__I0
timestamp 1669390400
transform 1 0 70560 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__S0
timestamp 1669390400
transform 1 0 70784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__S1
timestamp 1669390400
transform 1 0 70112 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A1
timestamp 1669390400
transform -1 0 70000 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0904__A2
timestamp 1669390400
transform 1 0 69216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__I
timestamp 1669390400
transform -1 0 67872 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__I
timestamp 1669390400
transform -1 0 65968 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__I1
timestamp 1669390400
transform 1 0 71120 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__I2
timestamp 1669390400
transform 1 0 70672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__S0
timestamp 1669390400
transform -1 0 71008 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__S1
timestamp 1669390400
transform 1 0 72016 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__I
timestamp 1669390400
transform -1 0 71232 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A1
timestamp 1669390400
transform 1 0 68544 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__B
timestamp 1669390400
transform 1 0 68096 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__I
timestamp 1669390400
transform 1 0 72464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0911__I
timestamp 1669390400
transform -1 0 70448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__I0
timestamp 1669390400
transform 1 0 74368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__I3
timestamp 1669390400
transform 1 0 74032 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__S0
timestamp 1669390400
transform 1 0 73472 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__S1
timestamp 1669390400
transform 1 0 73920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A1
timestamp 1669390400
transform -1 0 72016 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0913__A2
timestamp 1669390400
transform -1 0 71680 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__I
timestamp 1669390400
transform 1 0 68432 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__I1
timestamp 1669390400
transform 1 0 69328 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__I2
timestamp 1669390400
transform 1 0 69776 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__I3
timestamp 1669390400
transform 1 0 70224 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__S0
timestamp 1669390400
transform 1 0 69328 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0916__I
timestamp 1669390400
transform -1 0 70560 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0917__A1
timestamp 1669390400
transform 1 0 69216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__I1
timestamp 1669390400
transform 1 0 56672 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__S0
timestamp 1669390400
transform 1 0 61152 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__S1
timestamp 1669390400
transform 1 0 61600 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__A1
timestamp 1669390400
transform 1 0 59024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__A2
timestamp 1669390400
transform -1 0 58352 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__I2
timestamp 1669390400
transform 1 0 58912 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__S0
timestamp 1669390400
transform 1 0 61152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__S1
timestamp 1669390400
transform 1 0 61600 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__A1
timestamp 1669390400
transform 1 0 59248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__B
timestamp 1669390400
transform -1 0 59584 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__I0
timestamp 1669390400
transform 1 0 57344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__I1
timestamp 1669390400
transform -1 0 62720 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__I2
timestamp 1669390400
transform 1 0 62944 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__S0
timestamp 1669390400
transform 1 0 61600 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__S1
timestamp 1669390400
transform 1 0 62048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A1
timestamp 1669390400
transform 1 0 60256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A2
timestamp 1669390400
transform -1 0 60032 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__I0
timestamp 1669390400
transform -1 0 62272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__I1
timestamp 1669390400
transform 1 0 67200 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__I3
timestamp 1669390400
transform 1 0 66752 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__S0
timestamp 1669390400
transform 1 0 66304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__A1
timestamp 1669390400
transform 1 0 63952 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__I0
timestamp 1669390400
transform -1 0 62384 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__S0
timestamp 1669390400
transform 1 0 61264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__S1
timestamp 1669390400
transform 1 0 61712 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1669390400
transform 1 0 61712 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A2
timestamp 1669390400
transform 1 0 61264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__I
timestamp 1669390400
transform 1 0 81200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__I
timestamp 1669390400
transform -1 0 72800 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__I2
timestamp 1669390400
transform 1 0 54992 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__S0
timestamp 1669390400
transform 1 0 56672 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__S1
timestamp 1669390400
transform 1 0 58464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__A1
timestamp 1669390400
transform -1 0 58688 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0933__B
timestamp 1669390400
transform -1 0 58688 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__I1
timestamp 1669390400
transform 1 0 59696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__I2
timestamp 1669390400
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__S0
timestamp 1669390400
transform -1 0 59024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__S1
timestamp 1669390400
transform -1 0 59472 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A1
timestamp 1669390400
transform 1 0 60144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0935__A2
timestamp 1669390400
transform 1 0 59696 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__I0
timestamp 1669390400
transform 1 0 65744 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__I1
timestamp 1669390400
transform 1 0 66640 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__I3
timestamp 1669390400
transform 1 0 65968 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__S0
timestamp 1669390400
transform 1 0 65520 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__A1
timestamp 1669390400
transform 1 0 62944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__S0
timestamp 1669390400
transform 1 0 62944 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__S1
timestamp 1669390400
transform 1 0 63392 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A1
timestamp 1669390400
transform -1 0 58800 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A2
timestamp 1669390400
transform 1 0 59360 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__I1
timestamp 1669390400
transform 1 0 52864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__I2
timestamp 1669390400
transform 1 0 53312 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__S0
timestamp 1669390400
transform 1 0 56672 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__S1
timestamp 1669390400
transform -1 0 57568 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__A1
timestamp 1669390400
transform 1 0 59360 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__B
timestamp 1669390400
transform 1 0 59808 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__I0
timestamp 1669390400
transform -1 0 54432 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__I1
timestamp 1669390400
transform 1 0 53312 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__I2
timestamp 1669390400
transform 1 0 53760 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__S0
timestamp 1669390400
transform 1 0 58240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0943__S1
timestamp 1669390400
transform 1 0 58688 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__A1
timestamp 1669390400
transform 1 0 55664 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0944__A2
timestamp 1669390400
transform 1 0 56112 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__I0
timestamp 1669390400
transform -1 0 65968 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__I1
timestamp 1669390400
transform 1 0 66192 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0945__S0
timestamp 1669390400
transform 1 0 65296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0946__A1
timestamp 1669390400
transform 1 0 63392 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__I
timestamp 1669390400
transform -1 0 81760 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0949__I
timestamp 1669390400
transform 1 0 70784 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A1
timestamp 1669390400
transform 1 0 76272 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__I
timestamp 1669390400
transform 1 0 77168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A1
timestamp 1669390400
transform -1 0 71232 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__I
timestamp 1669390400
transform 1 0 77616 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__I0
timestamp 1669390400
transform 1 0 83888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__S
timestamp 1669390400
transform 1 0 80640 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0958__S
timestamp 1669390400
transform -1 0 79296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0960__I
timestamp 1669390400
transform 1 0 82544 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__I0
timestamp 1669390400
transform 1 0 85120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__S
timestamp 1669390400
transform 1 0 82320 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0963__S
timestamp 1669390400
transform 1 0 84448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0965__I
timestamp 1669390400
transform 1 0 81200 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__I
timestamp 1669390400
transform 1 0 68768 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__I0
timestamp 1669390400
transform 1 0 83664 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__S
timestamp 1669390400
transform -1 0 81536 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__S
timestamp 1669390400
transform 1 0 82880 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__I
timestamp 1669390400
transform -1 0 66192 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__I0
timestamp 1669390400
transform 1 0 67200 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0972__S
timestamp 1669390400
transform -1 0 67872 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__I0
timestamp 1669390400
transform 1 0 87024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__S
timestamp 1669390400
transform -1 0 84672 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__I
timestamp 1669390400
transform 1 0 47824 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__I
timestamp 1669390400
transform 1 0 67984 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0978__I0
timestamp 1669390400
transform -1 0 48944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0978__S
timestamp 1669390400
transform 1 0 51072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__S
timestamp 1669390400
transform 1 0 68544 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__I
timestamp 1669390400
transform 1 0 46928 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__I0
timestamp 1669390400
transform -1 0 48048 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__S
timestamp 1669390400
transform 1 0 51968 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__I0
timestamp 1669390400
transform 1 0 51408 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0985__S
timestamp 1669390400
transform 1 0 51856 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__I
timestamp 1669390400
transform 1 0 52528 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__I
timestamp 1669390400
transform -1 0 74816 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__I0
timestamp 1669390400
transform 1 0 51072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__S
timestamp 1669390400
transform 1 0 52192 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__S
timestamp 1669390400
transform 1 0 53872 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__I0
timestamp 1669390400
transform 1 0 52528 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0993__S
timestamp 1669390400
transform 1 0 53424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__I
timestamp 1669390400
transform 1 0 93296 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__I
timestamp 1669390400
transform 1 0 72016 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A1
timestamp 1669390400
transform 1 0 79296 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A2
timestamp 1669390400
transform 1 0 77392 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0997__A3
timestamp 1669390400
transform 1 0 68544 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__I
timestamp 1669390400
transform 1 0 76160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__I0
timestamp 1669390400
transform -1 0 93968 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__S
timestamp 1669390400
transform -1 0 93408 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__S
timestamp 1669390400
transform 1 0 77728 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__I
timestamp 1669390400
transform 1 0 89824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1004__S
timestamp 1669390400
transform 1 0 88704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__I0
timestamp 1669390400
transform 1 0 92400 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__S
timestamp 1669390400
transform 1 0 98000 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1008__I
timestamp 1669390400
transform 1 0 82432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__I
timestamp 1669390400
transform 1 0 73248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__I0
timestamp 1669390400
transform 1 0 84560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__S
timestamp 1669390400
transform -1 0 82656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__I0
timestamp 1669390400
transform 1 0 87472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__S
timestamp 1669390400
transform -1 0 85344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__I
timestamp 1669390400
transform 1 0 68992 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1015__I0
timestamp 1669390400
transform 1 0 71792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1015__S
timestamp 1669390400
transform 1 0 71344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__I0
timestamp 1669390400
transform 1 0 85120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__S
timestamp 1669390400
transform 1 0 82656 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__I
timestamp 1669390400
transform 1 0 57344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1020__I
timestamp 1669390400
transform 1 0 70784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__I0
timestamp 1669390400
transform 1 0 61488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__S
timestamp 1669390400
transform -1 0 65632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__I0
timestamp 1669390400
transform -1 0 68768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__S
timestamp 1669390400
transform 1 0 70336 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__I
timestamp 1669390400
transform 1 0 54208 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__I0
timestamp 1669390400
transform 1 0 58128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__S
timestamp 1669390400
transform 1 0 60256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__I0
timestamp 1669390400
transform 1 0 62496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1028__S
timestamp 1669390400
transform 1 0 65520 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__I
timestamp 1669390400
transform 1 0 50512 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__I
timestamp 1669390400
transform 1 0 71344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__I0
timestamp 1669390400
transform 1 0 53312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__S
timestamp 1669390400
transform 1 0 53760 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__I0
timestamp 1669390400
transform 1 0 59248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__S
timestamp 1669390400
transform 1 0 59248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__I
timestamp 1669390400
transform 1 0 75264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A1
timestamp 1669390400
transform 1 0 71120 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A2
timestamp 1669390400
transform 1 0 76496 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__I
timestamp 1669390400
transform -1 0 71120 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A1
timestamp 1669390400
transform 1 0 76160 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__I
timestamp 1669390400
transform 1 0 73696 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1669390400
transform 1 0 75040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A2
timestamp 1669390400
transform -1 0 73472 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A1
timestamp 1669390400
transform 1 0 76272 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A2
timestamp 1669390400
transform -1 0 73472 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__I
timestamp 1669390400
transform 1 0 73696 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A2
timestamp 1669390400
transform 1 0 76048 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__I0
timestamp 1669390400
transform -1 0 54432 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__S
timestamp 1669390400
transform -1 0 53536 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__I
timestamp 1669390400
transform 1 0 84000 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1669390400
transform -1 0 80416 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A3
timestamp 1669390400
transform -1 0 68320 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__I
timestamp 1669390400
transform 1 0 77392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I0
timestamp 1669390400
transform 1 0 96880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__S
timestamp 1669390400
transform 1 0 93184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__I0
timestamp 1669390400
transform -1 0 81424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__S
timestamp 1669390400
transform 1 0 78512 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__S
timestamp 1669390400
transform 1 0 88480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__I0
timestamp 1669390400
transform -1 0 93856 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__S
timestamp 1669390400
transform 1 0 97104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__I
timestamp 1669390400
transform 1 0 74592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__I0
timestamp 1669390400
transform 1 0 86016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__S
timestamp 1669390400
transform 1 0 88592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__I0
timestamp 1669390400
transform -1 0 90384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__S
timestamp 1669390400
transform 1 0 88480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__I0
timestamp 1669390400
transform 1 0 73024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__S
timestamp 1669390400
transform -1 0 75152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__I0
timestamp 1669390400
transform 1 0 87024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__S
timestamp 1669390400
transform 1 0 84896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__I
timestamp 1669390400
transform -1 0 73472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__I0
timestamp 1669390400
transform -1 0 61488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__S
timestamp 1669390400
transform -1 0 63616 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__I0
timestamp 1669390400
transform 1 0 73472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1072__S
timestamp 1669390400
transform 1 0 72576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__I0
timestamp 1669390400
transform 1 0 61488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__S
timestamp 1669390400
transform 1 0 63616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__I0
timestamp 1669390400
transform 1 0 64512 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__S
timestamp 1669390400
transform 1 0 66640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__I
timestamp 1669390400
transform 1 0 76384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__I0
timestamp 1669390400
transform 1 0 62720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__S
timestamp 1669390400
transform 1 0 65296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__I0
timestamp 1669390400
transform -1 0 65520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__S
timestamp 1669390400
transform -1 0 65072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__I0
timestamp 1669390400
transform -1 0 72800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__S
timestamp 1669390400
transform 1 0 69328 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__I0
timestamp 1669390400
transform 1 0 65744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__S
timestamp 1669390400
transform 1 0 65296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__I
timestamp 1669390400
transform 1 0 93520 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__A1
timestamp 1669390400
transform 1 0 77168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1669390400
transform 1 0 71680 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A2
timestamp 1669390400
transform -1 0 72016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A4
timestamp 1669390400
transform 1 0 77168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__I
timestamp 1669390400
transform 1 0 77616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A1
timestamp 1669390400
transform 1 0 95984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1092__A2
timestamp 1669390400
transform -1 0 95760 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__I
timestamp 1669390400
transform -1 0 70112 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A1
timestamp 1669390400
transform 1 0 73472 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A2
timestamp 1669390400
transform 1 0 72576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A4
timestamp 1669390400
transform -1 0 72352 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__A2
timestamp 1669390400
transform -1 0 96656 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1669390400
transform 1 0 82432 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A2
timestamp 1669390400
transform 1 0 81984 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A2
timestamp 1669390400
transform 1 0 78736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__I
timestamp 1669390400
transform 1 0 90832 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A1
timestamp 1669390400
transform -1 0 94416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A2
timestamp 1669390400
transform -1 0 94864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A2
timestamp 1669390400
transform 1 0 97216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A2
timestamp 1669390400
transform -1 0 95200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1105__I
timestamp 1669390400
transform 1 0 75264 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1669390400
transform 1 0 92624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A2
timestamp 1669390400
transform 1 0 93520 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__I
timestamp 1669390400
transform 1 0 89936 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__A2
timestamp 1669390400
transform 1 0 97888 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__A2
timestamp 1669390400
transform 1 0 97552 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__A2
timestamp 1669390400
transform -1 0 93296 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__A1
timestamp 1669390400
transform -1 0 93296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__I
timestamp 1669390400
transform 1 0 67648 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__I
timestamp 1669390400
transform 1 0 76832 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A2
timestamp 1669390400
transform -1 0 68992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A2
timestamp 1669390400
transform -1 0 72800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1669390400
transform 1 0 97104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A2
timestamp 1669390400
transform 1 0 93968 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__I
timestamp 1669390400
transform 1 0 58128 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__A1
timestamp 1669390400
transform 1 0 60592 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__A2
timestamp 1669390400
transform 1 0 66864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1124__A2
timestamp 1669390400
transform 1 0 66976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A2
timestamp 1669390400
transform 1 0 74480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__I
timestamp 1669390400
transform 1 0 55440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1669390400
transform 1 0 62048 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A2
timestamp 1669390400
transform -1 0 61376 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1130__A2
timestamp 1669390400
transform -1 0 66304 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__I
timestamp 1669390400
transform 1 0 77168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A1
timestamp 1669390400
transform 1 0 66864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A2
timestamp 1669390400
transform -1 0 67536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__I
timestamp 1669390400
transform 1 0 50960 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__A1
timestamp 1669390400
transform 1 0 60592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__A2
timestamp 1669390400
transform -1 0 61040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A2
timestamp 1669390400
transform 1 0 67312 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A1
timestamp 1669390400
transform 1 0 65296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A2
timestamp 1669390400
transform 1 0 64512 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__I
timestamp 1669390400
transform 1 0 77616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__I0
timestamp 1669390400
transform 1 0 77168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__S
timestamp 1669390400
transform 1 0 77840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__A1
timestamp 1669390400
transform 1 0 65968 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1144__A2
timestamp 1669390400
transform 1 0 66416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__I
timestamp 1669390400
transform 1 0 80192 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__A2
timestamp 1669390400
transform 1 0 77840 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A1
timestamp 1669390400
transform 1 0 94976 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A2
timestamp 1669390400
transform -1 0 94192 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__A2
timestamp 1669390400
transform 1 0 79744 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__I
timestamp 1669390400
transform 1 0 80640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__A2
timestamp 1669390400
transform 1 0 97328 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A2
timestamp 1669390400
transform -1 0 82656 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__A2
timestamp 1669390400
transform 1 0 81984 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__A1
timestamp 1669390400
transform 1 0 93072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__A2
timestamp 1669390400
transform -1 0 92400 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__A2
timestamp 1669390400
transform 1 0 96880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__A2
timestamp 1669390400
transform 1 0 97104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A2
timestamp 1669390400
transform -1 0 93744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A2
timestamp 1669390400
transform 1 0 96320 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A2
timestamp 1669390400
transform -1 0 93744 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A2
timestamp 1669390400
transform 1 0 66976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__I
timestamp 1669390400
transform 1 0 70112 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__A2
timestamp 1669390400
transform -1 0 68992 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__A2
timestamp 1669390400
transform -1 0 95760 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A1
timestamp 1669390400
transform -1 0 57232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A2
timestamp 1669390400
transform 1 0 57456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A2
timestamp 1669390400
transform 1 0 58912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A2
timestamp 1669390400
transform -1 0 70784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1181__A1
timestamp 1669390400
transform 1 0 57344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1181__A2
timestamp 1669390400
transform 1 0 57792 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A2
timestamp 1669390400
transform 1 0 59136 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__A2
timestamp 1669390400
transform 1 0 58912 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A1
timestamp 1669390400
transform 1 0 54992 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A2
timestamp 1669390400
transform 1 0 57008 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__A2
timestamp 1669390400
transform 1 0 58688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A2
timestamp 1669390400
transform 1 0 57792 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1192__I
timestamp 1669390400
transform 1 0 81872 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1669390400
transform 1 0 77616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A2
timestamp 1669390400
transform 1 0 77168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__A2
timestamp 1669390400
transform 1 0 57344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1197__I
timestamp 1669390400
transform 1 0 95200 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A1
timestamp 1669390400
transform 1 0 83216 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A3
timestamp 1669390400
transform -1 0 74592 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A4
timestamp 1669390400
transform 1 0 83664 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1200__I
timestamp 1669390400
transform -1 0 75824 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__I1
timestamp 1669390400
transform 1 0 97104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__S
timestamp 1669390400
transform 1 0 97104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__I1
timestamp 1669390400
transform -1 0 80080 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__S
timestamp 1669390400
transform -1 0 77952 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1205__I
timestamp 1669390400
transform -1 0 92624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__I1
timestamp 1669390400
transform 1 0 96320 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__S
timestamp 1669390400
transform 1 0 93968 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1208__I1
timestamp 1669390400
transform -1 0 94304 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1208__S
timestamp 1669390400
transform 1 0 93632 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__I
timestamp 1669390400
transform 1 0 87136 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__I
timestamp 1669390400
transform 1 0 73696 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__I1
timestamp 1669390400
transform 1 0 92064 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__S
timestamp 1669390400
transform -1 0 89152 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__I1
timestamp 1669390400
transform 1 0 93520 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__S
timestamp 1669390400
transform 1 0 93072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__I
timestamp 1669390400
transform -1 0 68096 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__I1
timestamp 1669390400
transform 1 0 70112 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__S
timestamp 1669390400
transform 1 0 72240 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__I1
timestamp 1669390400
transform -1 0 91392 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__S
timestamp 1669390400
transform 1 0 91056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__I
timestamp 1669390400
transform -1 0 53424 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__I
timestamp 1669390400
transform 1 0 72464 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__I1
timestamp 1669390400
transform 1 0 57792 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__S
timestamp 1669390400
transform 1 0 59472 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__I1
timestamp 1669390400
transform 1 0 71120 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1225__S
timestamp 1669390400
transform -1 0 71344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__I
timestamp 1669390400
transform 1 0 54768 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__I1
timestamp 1669390400
transform -1 0 54768 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__S
timestamp 1669390400
transform 1 0 58240 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__S
timestamp 1669390400
transform 1 0 59696 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__I
timestamp 1669390400
transform -1 0 51744 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__I
timestamp 1669390400
transform 1 0 76608 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1234__I1
timestamp 1669390400
transform 1 0 53088 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1234__S
timestamp 1669390400
transform -1 0 53760 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__S
timestamp 1669390400
transform 1 0 59696 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A1
timestamp 1669390400
transform 1 0 81088 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1238__A2
timestamp 1669390400
transform 1 0 81536 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__I1
timestamp 1669390400
transform -1 0 52752 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1240__S
timestamp 1669390400
transform 1 0 52080 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A1
timestamp 1669390400
transform 1 0 81648 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A2
timestamp 1669390400
transform 1 0 78848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A3
timestamp 1669390400
transform 1 0 79744 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1242__A4
timestamp 1669390400
transform 1 0 82096 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__I
timestamp 1669390400
transform 1 0 76496 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__I1
timestamp 1669390400
transform 1 0 94976 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1244__S
timestamp 1669390400
transform -1 0 94752 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__I1
timestamp 1669390400
transform -1 0 79744 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__S
timestamp 1669390400
transform -1 0 78736 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__I1
timestamp 1669390400
transform -1 0 94528 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1248__S
timestamp 1669390400
transform 1 0 94304 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1250__I1
timestamp 1669390400
transform -1 0 97328 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1250__S
timestamp 1669390400
transform 1 0 94304 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__I
timestamp 1669390400
transform -1 0 72800 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1253__I1
timestamp 1669390400
transform 1 0 90944 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1253__S
timestamp 1669390400
transform 1 0 90496 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__I1
timestamp 1669390400
transform 1 0 97776 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__S
timestamp 1669390400
transform 1 0 96880 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__I1
timestamp 1669390400
transform -1 0 71120 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__S
timestamp 1669390400
transform 1 0 73696 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1259__S
timestamp 1669390400
transform 1 0 90496 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1261__I
timestamp 1669390400
transform -1 0 75152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__I1
timestamp 1669390400
transform -1 0 57568 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__S
timestamp 1669390400
transform -1 0 59696 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__I1
timestamp 1669390400
transform 1 0 71680 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__S
timestamp 1669390400
transform 1 0 73248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__I1
timestamp 1669390400
transform 1 0 60592 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__S
timestamp 1669390400
transform -1 0 64512 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__S
timestamp 1669390400
transform 1 0 60256 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__I
timestamp 1669390400
transform -1 0 75600 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__I1
timestamp 1669390400
transform 1 0 65744 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__S
timestamp 1669390400
transform 1 0 67648 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__I1
timestamp 1669390400
transform -1 0 63168 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__S
timestamp 1669390400
transform 1 0 65296 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__I
timestamp 1669390400
transform -1 0 76384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__I1
timestamp 1669390400
transform 1 0 77168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__S
timestamp 1669390400
transform 1 0 76496 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1278__S
timestamp 1669390400
transform 1 0 65072 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1669390400
transform -1 0 78736 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A2
timestamp 1669390400
transform 1 0 75712 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__I
timestamp 1669390400
transform 1 0 74256 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__I1
timestamp 1669390400
transform -1 0 94752 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__S
timestamp 1669390400
transform 1 0 92176 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__S
timestamp 1669390400
transform -1 0 79296 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__I1
timestamp 1669390400
transform 1 0 97328 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__S
timestamp 1669390400
transform 1 0 92400 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__S
timestamp 1669390400
transform 1 0 93520 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__I
timestamp 1669390400
transform 1 0 73584 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__I1
timestamp 1669390400
transform 1 0 89264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__S
timestamp 1669390400
transform -1 0 87136 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__S
timestamp 1669390400
transform 1 0 87584 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__I1
timestamp 1669390400
transform 1 0 69888 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__S
timestamp 1669390400
transform 1 0 71568 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1297__S
timestamp 1669390400
transform 1 0 89152 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__I
timestamp 1669390400
transform -1 0 72912 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__I1
timestamp 1669390400
transform -1 0 56112 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__S
timestamp 1669390400
transform -1 0 54880 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__S
timestamp 1669390400
transform 1 0 70672 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1304__I1
timestamp 1669390400
transform 1 0 57344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1304__S
timestamp 1669390400
transform 1 0 57680 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__I1
timestamp 1669390400
transform -1 0 55664 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__S
timestamp 1669390400
transform 1 0 54992 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__I
timestamp 1669390400
transform 1 0 73808 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__I1
timestamp 1669390400
transform 1 0 62608 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__S
timestamp 1669390400
transform -1 0 64400 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1311__S
timestamp 1669390400
transform 1 0 60256 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__I1
timestamp 1669390400
transform -1 0 76608 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__S
timestamp 1669390400
transform 1 0 74480 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__S
timestamp 1669390400
transform 1 0 64400 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A2
timestamp 1669390400
transform 1 0 72800 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__I
timestamp 1669390400
transform 1 0 76272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__I0
timestamp 1669390400
transform 1 0 98000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__I1
timestamp 1669390400
transform 1 0 96096 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1320__S
timestamp 1669390400
transform 1 0 97104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__I0
timestamp 1669390400
transform -1 0 77168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1322__S
timestamp 1669390400
transform 1 0 76496 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__I1
timestamp 1669390400
transform -1 0 89824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1324__S
timestamp 1669390400
transform 1 0 90048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__I0
timestamp 1669390400
transform 1 0 93968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__I1
timestamp 1669390400
transform 1 0 93520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1326__S
timestamp 1669390400
transform -1 0 90720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__I
timestamp 1669390400
transform 1 0 72240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__I0
timestamp 1669390400
transform 1 0 84336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1329__S
timestamp 1669390400
transform -1 0 80752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__I0
timestamp 1669390400
transform 1 0 84224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__I1
timestamp 1669390400
transform 1 0 83776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1331__S
timestamp 1669390400
transform -1 0 81648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__I0
timestamp 1669390400
transform 1 0 71568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__S
timestamp 1669390400
transform 1 0 71120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__I0
timestamp 1669390400
transform 1 0 81648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__S
timestamp 1669390400
transform 1 0 81200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__I
timestamp 1669390400
transform 1 0 70672 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__I0
timestamp 1669390400
transform 1 0 61040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1338__S
timestamp 1669390400
transform -1 0 59808 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__I0
timestamp 1669390400
transform 1 0 69664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__S
timestamp 1669390400
transform 1 0 69216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__I0
timestamp 1669390400
transform 1 0 55664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__S
timestamp 1669390400
transform 1 0 58016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__I0
timestamp 1669390400
transform 1 0 59808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__S
timestamp 1669390400
transform 1 0 59360 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__I
timestamp 1669390400
transform 1 0 72688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__I0
timestamp 1669390400
transform 1 0 54656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__S
timestamp 1669390400
transform 1 0 54208 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__I0
timestamp 1669390400
transform -1 0 56672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__S
timestamp 1669390400
transform 1 0 56896 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__I1
timestamp 1669390400
transform 1 0 74816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__S
timestamp 1669390400
transform 1 0 73808 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__I0
timestamp 1669390400
transform 1 0 54768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__S
timestamp 1669390400
transform 1 0 55104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1355__I
timestamp 1669390400
transform -1 0 81648 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A3
timestamp 1669390400
transform -1 0 75488 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__I
timestamp 1669390400
transform 1 0 76160 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A1
timestamp 1669390400
transform -1 0 94192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__A2
timestamp 1669390400
transform 1 0 96768 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__I
timestamp 1669390400
transform 1 0 82320 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A1
timestamp 1669390400
transform 1 0 82656 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A3
timestamp 1669390400
transform 1 0 82208 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__A4
timestamp 1669390400
transform -1 0 75488 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__I
timestamp 1669390400
transform -1 0 76496 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__A2
timestamp 1669390400
transform 1 0 91280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A2
timestamp 1669390400
transform -1 0 78064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__A2
timestamp 1669390400
transform -1 0 75152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A1
timestamp 1669390400
transform 1 0 91840 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A2
timestamp 1669390400
transform -1 0 92512 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A2
timestamp 1669390400
transform -1 0 92512 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__I
timestamp 1669390400
transform 1 0 71008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__A2
timestamp 1669390400
transform -1 0 87360 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A2
timestamp 1669390400
transform 1 0 89264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A2
timestamp 1669390400
transform 1 0 92400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1669390400
transform -1 0 89040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A1
timestamp 1669390400
transform 1 0 86240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__A2
timestamp 1669390400
transform -1 0 85904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__I
timestamp 1669390400
transform 1 0 70448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__A2
timestamp 1669390400
transform 1 0 67760 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1382__I
timestamp 1669390400
transform 1 0 77168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1383__A2
timestamp 1669390400
transform 1 0 71232 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A2
timestamp 1669390400
transform 1 0 84336 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A1
timestamp 1669390400
transform -1 0 83552 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__A1
timestamp 1669390400
transform -1 0 57568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1387__A2
timestamp 1669390400
transform 1 0 59696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1388__A2
timestamp 1669390400
transform 1 0 59472 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A1
timestamp 1669390400
transform 1 0 70112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A2
timestamp 1669390400
transform 1 0 70784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A1
timestamp 1669390400
transform 1 0 56000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__A2
timestamp 1669390400
transform -1 0 55776 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1393__A2
timestamp 1669390400
transform -1 0 54320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1395__I
timestamp 1669390400
transform 1 0 71680 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A2
timestamp 1669390400
transform 1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A1
timestamp 1669390400
transform 1 0 53088 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A2
timestamp 1669390400
transform -1 0 54880 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A2
timestamp 1669390400
transform -1 0 55328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A2
timestamp 1669390400
transform -1 0 55328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__I0
timestamp 1669390400
transform 1 0 74592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__S
timestamp 1669390400
transform 1 0 74144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__A2
timestamp 1669390400
transform -1 0 54880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1407__A1
timestamp 1669390400
transform -1 0 72576 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1407__A3
timestamp 1669390400
transform -1 0 72128 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__I
timestamp 1669390400
transform -1 0 75936 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1669390400
transform 1 0 91616 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A2
timestamp 1669390400
transform 1 0 86800 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1410__A3
timestamp 1669390400
transform 1 0 71568 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1410__A4
timestamp 1669390400
transform 1 0 71680 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__I
timestamp 1669390400
transform 1 0 77840 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A2
timestamp 1669390400
transform 1 0 92288 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__A2
timestamp 1669390400
transform -1 0 79632 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1669390400
transform -1 0 79184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A1
timestamp 1669390400
transform 1 0 92064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A2
timestamp 1669390400
transform -1 0 90608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A2
timestamp 1669390400
transform -1 0 90160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__I
timestamp 1669390400
transform 1 0 71120 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__A2
timestamp 1669390400
transform -1 0 86912 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A2
timestamp 1669390400
transform 1 0 91616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__A2
timestamp 1669390400
transform -1 0 93296 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1426__A2
timestamp 1669390400
transform 1 0 86352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__I
timestamp 1669390400
transform 1 0 69888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1429__A2
timestamp 1669390400
transform 1 0 68432 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__I
timestamp 1669390400
transform -1 0 71568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1669390400
transform 1 0 70784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A2
timestamp 1669390400
transform 1 0 87920 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A1
timestamp 1669390400
transform 1 0 62160 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A2
timestamp 1669390400
transform 1 0 63952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1436__A2
timestamp 1669390400
transform 1 0 66080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A2
timestamp 1669390400
transform 1 0 71232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A1
timestamp 1669390400
transform 1 0 59248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A2
timestamp 1669390400
transform 1 0 60256 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1669390400
transform 1 0 66080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1443__I
timestamp 1669390400
transform 1 0 76384 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__A2
timestamp 1669390400
transform -1 0 66528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__A1
timestamp 1669390400
transform 1 0 61152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__A2
timestamp 1669390400
transform 1 0 62608 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1447__A2
timestamp 1669390400
transform -1 0 64624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A2
timestamp 1669390400
transform 1 0 61264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__A2
timestamp 1669390400
transform -1 0 66976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__I0
timestamp 1669390400
transform 1 0 77280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__S
timestamp 1669390400
transform -1 0 74704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1453__A2
timestamp 1669390400
transform 1 0 66080 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A1
timestamp 1669390400
transform -1 0 61824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__A1
timestamp 1669390400
transform -1 0 72800 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__A2
timestamp 1669390400
transform 1 0 78848 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1455__A3
timestamp 1669390400
transform 1 0 80192 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__I
timestamp 1669390400
transform 1 0 77168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__I1
timestamp 1669390400
transform 1 0 93632 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__S
timestamp 1669390400
transform -1 0 96208 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__I1
timestamp 1669390400
transform 1 0 79968 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__S
timestamp 1669390400
transform -1 0 77840 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__I1
timestamp 1669390400
transform 1 0 97104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1461__S
timestamp 1669390400
transform 1 0 97552 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__I1
timestamp 1669390400
transform -1 0 93856 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__S
timestamp 1669390400
transform 1 0 94080 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__I
timestamp 1669390400
transform 1 0 74816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__I1
timestamp 1669390400
transform 1 0 93072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__S
timestamp 1669390400
transform -1 0 93744 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__I1
timestamp 1669390400
transform 1 0 97104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__S
timestamp 1669390400
transform 1 0 96432 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__I1
timestamp 1669390400
transform 1 0 71456 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__S
timestamp 1669390400
transform -1 0 76160 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__I1
timestamp 1669390400
transform 1 0 92064 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__S
timestamp 1669390400
transform 1 0 88032 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__I
timestamp 1669390400
transform -1 0 73472 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__I1
timestamp 1669390400
transform 1 0 59696 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__S
timestamp 1669390400
transform -1 0 64064 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__I1
timestamp 1669390400
transform -1 0 72912 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__S
timestamp 1669390400
transform 1 0 73248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__I1
timestamp 1669390400
transform 1 0 60816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__S
timestamp 1669390400
transform 1 0 63616 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__I1
timestamp 1669390400
transform 1 0 65744 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__S
timestamp 1669390400
transform 1 0 65296 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__I
timestamp 1669390400
transform 1 0 75264 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__I1
timestamp 1669390400
transform 1 0 63168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__S
timestamp 1669390400
transform 1 0 63504 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__I1
timestamp 1669390400
transform 1 0 64288 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__S
timestamp 1669390400
transform 1 0 63840 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A1
timestamp 1669390400
transform 1 0 77616 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1669390400
transform 1 0 79408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__S
timestamp 1669390400
transform 1 0 63280 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A1
timestamp 1669390400
transform 1 0 70896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__I
timestamp 1669390400
transform -1 0 75600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__I0
timestamp 1669390400
transform -1 0 94752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__S
timestamp 1669390400
transform 1 0 94080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__I0
timestamp 1669390400
transform -1 0 76272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__S
timestamp 1669390400
transform -1 0 76496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__S
timestamp 1669390400
transform -1 0 89936 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__I0
timestamp 1669390400
transform 1 0 97104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__S
timestamp 1669390400
transform 1 0 93632 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__I
timestamp 1669390400
transform -1 0 74368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__I0
timestamp 1669390400
transform -1 0 83776 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__S
timestamp 1669390400
transform -1 0 83328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I0
timestamp 1669390400
transform -1 0 89376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__S
timestamp 1669390400
transform 1 0 91504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__I0
timestamp 1669390400
transform -1 0 70448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__S
timestamp 1669390400
transform 1 0 71344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__I0
timestamp 1669390400
transform -1 0 88592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1509__S
timestamp 1669390400
transform 1 0 85568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__I
timestamp 1669390400
transform -1 0 73920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__I0
timestamp 1669390400
transform 1 0 59696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__S
timestamp 1669390400
transform 1 0 59696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__I0
timestamp 1669390400
transform 1 0 69664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__S
timestamp 1669390400
transform -1 0 69440 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__I0
timestamp 1669390400
transform -1 0 53872 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__S
timestamp 1669390400
transform 1 0 53760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__I0
timestamp 1669390400
transform -1 0 58016 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1518__S
timestamp 1669390400
transform -1 0 57120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__I
timestamp 1669390400
transform 1 0 74144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__I0
timestamp 1669390400
transform 1 0 53760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__S
timestamp 1669390400
transform 1 0 53312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__I0
timestamp 1669390400
transform -1 0 53536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__S
timestamp 1669390400
transform 1 0 55216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__I1
timestamp 1669390400
transform 1 0 79072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__S
timestamp 1669390400
transform 1 0 75712 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__I0
timestamp 1669390400
transform -1 0 53536 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__S
timestamp 1669390400
transform 1 0 52976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A3
timestamp 1669390400
transform -1 0 74032 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A1
timestamp 1669390400
transform 1 0 83776 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A1
timestamp 1669390400
transform 1 0 83888 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A3
timestamp 1669390400
transform 1 0 80304 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__A4
timestamp 1669390400
transform 1 0 81872 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A2
timestamp 1669390400
transform 1 0 84672 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A2
timestamp 1669390400
transform 1 0 79520 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__A1
timestamp 1669390400
transform 1 0 84224 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__A2
timestamp 1669390400
transform 1 0 84224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A2
timestamp 1669390400
transform -1 0 90944 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__A1
timestamp 1669390400
transform 1 0 82656 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A2
timestamp 1669390400
transform -1 0 87808 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__A2
timestamp 1669390400
transform 1 0 91392 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1669390400
transform 1 0 69216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1669390400
transform 1 0 69888 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__A2
timestamp 1669390400
transform -1 0 69664 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1669390400
transform -1 0 91392 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A1
timestamp 1669390400
transform 1 0 52640 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A2
timestamp 1669390400
transform 1 0 53760 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1558__A2
timestamp 1669390400
transform 1 0 54208 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__A2
timestamp 1669390400
transform -1 0 70672 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1669390400
transform 1 0 48272 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A2
timestamp 1669390400
transform -1 0 48944 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A2
timestamp 1669390400
transform -1 0 49840 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A2
timestamp 1669390400
transform 1 0 55776 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A1
timestamp 1669390400
transform 1 0 52192 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__A2
timestamp 1669390400
transform 1 0 53312 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__A2
timestamp 1669390400
transform 1 0 53760 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A2
timestamp 1669390400
transform 1 0 54544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__I0
timestamp 1669390400
transform 1 0 77280 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__S
timestamp 1669390400
transform -1 0 75376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__A2
timestamp 1669390400
transform 1 0 55440 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A1
timestamp 1669390400
transform 1 0 70560 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A3
timestamp 1669390400
transform 1 0 71344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A4
timestamp 1669390400
transform 1 0 76272 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__I
timestamp 1669390400
transform 1 0 75712 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1669390400
transform -1 0 82320 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A2
timestamp 1669390400
transform 1 0 83664 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A3
timestamp 1669390400
transform -1 0 75040 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A4
timestamp 1669390400
transform -1 0 66304 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__I
timestamp 1669390400
transform 1 0 72576 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A2
timestamp 1669390400
transform 1 0 80528 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A2
timestamp 1669390400
transform 1 0 76720 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A2
timestamp 1669390400
transform 1 0 75040 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A1
timestamp 1669390400
transform -1 0 84448 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A2
timestamp 1669390400
transform -1 0 84448 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1669390400
transform 1 0 83104 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I
timestamp 1669390400
transform -1 0 72128 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__A2
timestamp 1669390400
transform 1 0 80080 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1593__A1
timestamp 1669390400
transform 1 0 85120 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1593__A2
timestamp 1669390400
transform 1 0 84560 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A2
timestamp 1669390400
transform -1 0 81312 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__A2
timestamp 1669390400
transform -1 0 81536 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__I
timestamp 1669390400
transform 1 0 70560 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A1
timestamp 1669390400
transform -1 0 68656 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A2
timestamp 1669390400
transform 1 0 69216 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__I
timestamp 1669390400
transform 1 0 73248 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A2
timestamp 1669390400
transform 1 0 69776 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__A2
timestamp 1669390400
transform 1 0 80640 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1669390400
transform -1 0 49392 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A2
timestamp 1669390400
transform -1 0 49840 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A2
timestamp 1669390400
transform -1 0 53760 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__A2
timestamp 1669390400
transform 1 0 71456 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1669390400
transform 1 0 48272 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A2
timestamp 1669390400
transform -1 0 48944 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A2
timestamp 1669390400
transform 1 0 54544 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__I
timestamp 1669390400
transform -1 0 71232 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A2
timestamp 1669390400
transform 1 0 57568 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1669390400
transform 1 0 52640 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A2
timestamp 1669390400
transform -1 0 50288 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A2
timestamp 1669390400
transform -1 0 54544 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__A2
timestamp 1669390400
transform 1 0 55888 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A1
timestamp 1669390400
transform 1 0 81984 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A2
timestamp 1669390400
transform 1 0 76384 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A2
timestamp 1669390400
transform 1 0 57344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A1
timestamp 1669390400
transform 1 0 83776 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A2
timestamp 1669390400
transform -1 0 82768 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A2
timestamp 1669390400
transform -1 0 84448 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__I
timestamp 1669390400
transform -1 0 74368 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__A2
timestamp 1669390400
transform 1 0 77728 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1669390400
transform 1 0 84672 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A2
timestamp 1669390400
transform 1 0 84672 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1669390400
transform 1 0 85120 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A2
timestamp 1669390400
transform 1 0 86688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A1
timestamp 1669390400
transform -1 0 82320 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A2
timestamp 1669390400
transform 1 0 82768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1637__A2
timestamp 1669390400
transform 1 0 80528 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__A2
timestamp 1669390400
transform -1 0 85344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1669390400
transform 1 0 66192 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A1
timestamp 1669390400
transform -1 0 63616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A2
timestamp 1669390400
transform 1 0 63840 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1669390400
transform 1 0 72688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1669390400
transform 1 0 67984 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1669390400
transform 1 0 85568 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A1
timestamp 1669390400
transform 1 0 51856 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A2
timestamp 1669390400
transform 1 0 53312 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A2
timestamp 1669390400
transform -1 0 54880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1669390400
transform 1 0 67088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A2
timestamp 1669390400
transform 1 0 66864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A1
timestamp 1669390400
transform 1 0 50848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A2
timestamp 1669390400
transform 1 0 53088 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A2
timestamp 1669390400
transform -1 0 54432 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A2
timestamp 1669390400
transform 1 0 57344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A1
timestamp 1669390400
transform 1 0 51296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A2
timestamp 1669390400
transform -1 0 50288 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1660__A2
timestamp 1669390400
transform 1 0 56448 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A2
timestamp 1669390400
transform -1 0 54320 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1669390400
transform 1 0 58912 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A1
timestamp 1669390400
transform 1 0 72576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A2
timestamp 1669390400
transform 1 0 70784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__A2
timestamp 1669390400
transform 1 0 58576 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__A1
timestamp 1669390400
transform 1 0 58128 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A1
timestamp 1669390400
transform 1 0 73248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1669390400
transform -1 0 72016 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__CLK
timestamp 1669390400
transform 1 0 86016 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__CLK
timestamp 1669390400
transform 1 0 88144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__CLK
timestamp 1669390400
transform 1 0 80304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__CLK
timestamp 1669390400
transform 1 0 85120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__CLK
timestamp 1669390400
transform -1 0 51856 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__CLK
timestamp 1669390400
transform 1 0 51632 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__CLK
timestamp 1669390400
transform -1 0 53088 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__CLK
timestamp 1669390400
transform 1 0 50624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__CLK
timestamp 1669390400
transform 1 0 52080 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__CLK
timestamp 1669390400
transform 1 0 52864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__CLK
timestamp 1669390400
transform 1 0 94304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__CLK
timestamp 1669390400
transform -1 0 95648 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__CLK
timestamp 1669390400
transform 1 0 85120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__CLK
timestamp 1669390400
transform 1 0 88144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__CLK
timestamp 1669390400
transform 1 0 70672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__CLK
timestamp 1669390400
transform 1 0 85792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__CLK
timestamp 1669390400
transform 1 0 61264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__CLK
timestamp 1669390400
transform 1 0 61264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__CLK
timestamp 1669390400
transform 1 0 62160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__CLK
timestamp 1669390400
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__CLK
timestamp 1669390400
transform 1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__CLK
timestamp 1669390400
transform 1 0 76944 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__CLK
timestamp 1669390400
transform -1 0 53536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__CLK
timestamp 1669390400
transform 1 0 98000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__CLK
timestamp 1669390400
transform 1 0 77840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__CLK
timestamp 1669390400
transform 1 0 94528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__CLK
timestamp 1669390400
transform 1 0 73248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__CLK
timestamp 1669390400
transform 1 0 84448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__CLK
timestamp 1669390400
transform -1 0 60816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__CLK
timestamp 1669390400
transform -1 0 70672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__CLK
timestamp 1669390400
transform 1 0 64512 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__CLK
timestamp 1669390400
transform 1 0 66192 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__CLK
timestamp 1669390400
transform 1 0 65968 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__CLK
timestamp 1669390400
transform 1 0 65744 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__CLK
timestamp 1669390400
transform 1 0 72800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__CLK
timestamp 1669390400
transform 1 0 66416 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__CLK
timestamp 1669390400
transform -1 0 94752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__CLK
timestamp 1669390400
transform -1 0 82320 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__CLK
timestamp 1669390400
transform 1 0 97888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__CLK
timestamp 1669390400
transform -1 0 98112 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__CLK
timestamp 1669390400
transform 1 0 94752 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__CLK
timestamp 1669390400
transform 1 0 95088 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__CLK
timestamp 1669390400
transform 1 0 73248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__CLK
timestamp 1669390400
transform 1 0 98000 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__CLK
timestamp 1669390400
transform -1 0 75152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__CLK
timestamp 1669390400
transform 1 0 78960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__CLK
timestamp 1669390400
transform 1 0 96880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__CLK
timestamp 1669390400
transform -1 0 83104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__CLK
timestamp 1669390400
transform 1 0 97552 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__CLK
timestamp 1669390400
transform 1 0 97888 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__CLK
timestamp 1669390400
transform 1 0 65744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__CLK
timestamp 1669390400
transform 1 0 53424 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__CLK
timestamp 1669390400
transform 1 0 54320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__CLK
timestamp 1669390400
transform 1 0 58464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__CLK
timestamp 1669390400
transform 1 0 52640 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__CLK
timestamp 1669390400
transform 1 0 52640 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__CLK
timestamp 1669390400
transform 1 0 82320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__CLK
timestamp 1669390400
transform -1 0 52864 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__CLK
timestamp 1669390400
transform 1 0 80752 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__CLK
timestamp 1669390400
transform -1 0 94752 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__CLK
timestamp 1669390400
transform 1 0 91616 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__CLK
timestamp 1669390400
transform -1 0 92624 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__CLK
timestamp 1669390400
transform 1 0 71232 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__CLK
timestamp 1669390400
transform 1 0 93968 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__CLK
timestamp 1669390400
transform 1 0 60256 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__CLK
timestamp 1669390400
transform 1 0 70560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__CLK
timestamp 1669390400
transform -1 0 57568 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__CLK
timestamp 1669390400
transform 1 0 60368 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__CLK
timestamp 1669390400
transform 1 0 52080 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__CLK
timestamp 1669390400
transform 1 0 57344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__CLK
timestamp 1669390400
transform -1 0 82208 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__CLK
timestamp 1669390400
transform 1 0 52640 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__CLK
timestamp 1669390400
transform 1 0 80416 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__CLK
timestamp 1669390400
transform 1 0 73136 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__CLK
timestamp 1669390400
transform 1 0 60592 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__CLK
timestamp 1669390400
transform 1 0 70448 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__CLK
timestamp 1669390400
transform -1 0 63616 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__CLK
timestamp 1669390400
transform 1 0 62160 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__CLK
timestamp 1669390400
transform 1 0 66640 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__CLK
timestamp 1669390400
transform 1 0 64288 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__CLK
timestamp 1669390400
transform 1 0 77392 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__CLK
timestamp 1669390400
transform 1 0 65408 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__CLK
timestamp 1669390400
transform 1 0 78736 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__CLK
timestamp 1669390400
transform -1 0 90272 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__CLK
timestamp 1669390400
transform -1 0 71680 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__CLK
timestamp 1669390400
transform 1 0 90496 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__CLK
timestamp 1669390400
transform 1 0 54768 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__CLK
timestamp 1669390400
transform 1 0 69440 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__CLK
timestamp 1669390400
transform 1 0 53760 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__CLK
timestamp 1669390400
transform -1 0 54656 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__CLK
timestamp 1669390400
transform 1 0 64736 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__CLK
timestamp 1669390400
transform 1 0 60816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__CLK
timestamp 1669390400
transform 1 0 79744 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__CLK
timestamp 1669390400
transform 1 0 63952 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__CLK
timestamp 1669390400
transform 1 0 94192 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__CLK
timestamp 1669390400
transform 1 0 78176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__CLK
timestamp 1669390400
transform 1 0 97552 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__CLK
timestamp 1669390400
transform -1 0 70224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__CLK
timestamp 1669390400
transform 1 0 61040 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__CLK
timestamp 1669390400
transform 1 0 65296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__CLK
timestamp 1669390400
transform 1 0 53424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__CLK
timestamp 1669390400
transform 1 0 60256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__CLK
timestamp 1669390400
transform 1 0 53760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__CLK
timestamp 1669390400
transform 1 0 56672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__CLK
timestamp 1669390400
transform -1 0 77392 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__CLK
timestamp 1669390400
transform 1 0 53312 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__CLK
timestamp 1669390400
transform 1 0 93072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__CLK
timestamp 1669390400
transform -1 0 78736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__CLK
timestamp 1669390400
transform 1 0 91952 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__CLK
timestamp 1669390400
transform 1 0 93072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__CLK
timestamp 1669390400
transform -1 0 70224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__CLK
timestamp 1669390400
transform 1 0 84448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__CLK
timestamp 1669390400
transform 1 0 58688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__CLK
timestamp 1669390400
transform 1 0 70560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__CLK
timestamp 1669390400
transform 1 0 52864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__CLK
timestamp 1669390400
transform 1 0 56000 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__CLK
timestamp 1669390400
transform 1 0 52416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__CLK
timestamp 1669390400
transform -1 0 55776 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__CLK
timestamp 1669390400
transform 1 0 77168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__CLK
timestamp 1669390400
transform 1 0 52640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__CLK
timestamp 1669390400
transform 1 0 92400 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__CLK
timestamp 1669390400
transform -1 0 81424 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__CLK
timestamp 1669390400
transform 1 0 91168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__CLK
timestamp 1669390400
transform 1 0 91952 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__CLK
timestamp 1669390400
transform -1 0 92288 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__CLK
timestamp 1669390400
transform -1 0 66416 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__CLK
timestamp 1669390400
transform -1 0 91840 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__CLK
timestamp 1669390400
transform 1 0 64736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__CLK
timestamp 1669390400
transform -1 0 70784 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__CLK
timestamp 1669390400
transform 1 0 64736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__CLK
timestamp 1669390400
transform 1 0 65184 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__CLK
timestamp 1669390400
transform 1 0 65296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__CLK
timestamp 1669390400
transform -1 0 64624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__CLK
timestamp 1669390400
transform -1 0 77392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__CLK
timestamp 1669390400
transform 1 0 59808 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__CLK
timestamp 1669390400
transform 1 0 98000 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__CLK
timestamp 1669390400
transform 1 0 81200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__CLK
timestamp 1669390400
transform 1 0 96432 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__CLK
timestamp 1669390400
transform -1 0 97776 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__CLK
timestamp 1669390400
transform 1 0 94080 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__CLK
timestamp 1669390400
transform 1 0 97328 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__CLK
timestamp 1669390400
transform -1 0 94192 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__CLK
timestamp 1669390400
transform 1 0 64288 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__CLK
timestamp 1669390400
transform 1 0 64736 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__CLK
timestamp 1669390400
transform 1 0 65296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__CLK
timestamp 1669390400
transform 1 0 63056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__CLK
timestamp 1669390400
transform 1 0 63840 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__CLK
timestamp 1669390400
transform 1 0 80640 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__CLK
timestamp 1669390400
transform 1 0 63280 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__CLK
timestamp 1669390400
transform 1 0 68544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__CLK
timestamp 1669390400
transform 1 0 89152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__CLK
timestamp 1669390400
transform -1 0 58464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__CLK
timestamp 1669390400
transform 1 0 70896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__CLK
timestamp 1669390400
transform -1 0 53536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__CLK
timestamp 1669390400
transform 1 0 56672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__CLK
timestamp 1669390400
transform 1 0 52864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__CLK
timestamp 1669390400
transform 1 0 53760 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__CLK
timestamp 1669390400
transform 1 0 53760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__CLK
timestamp 1669390400
transform 1 0 65520 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__CLK
timestamp 1669390400
transform 1 0 52640 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__CLK
timestamp 1669390400
transform 1 0 54096 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__CLK
timestamp 1669390400
transform -1 0 57120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1889__CLK
timestamp 1669390400
transform -1 0 53536 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__CLK
timestamp 1669390400
transform 1 0 54544 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__CLK
timestamp 1669390400
transform -1 0 77392 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__CLK
timestamp 1669390400
transform 1 0 52640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__CLK
timestamp 1669390400
transform -1 0 82096 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__CLK
timestamp 1669390400
transform 1 0 77168 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__CLK
timestamp 1669390400
transform 1 0 79520 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__CLK
timestamp 1669390400
transform 1 0 85232 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__CLK
timestamp 1669390400
transform -1 0 84896 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__CLK
timestamp 1669390400
transform 1 0 86576 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__CLK
timestamp 1669390400
transform 1 0 69664 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__CLK
timestamp 1669390400
transform 1 0 82992 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__CLK
timestamp 1669390400
transform 1 0 53312 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__CLK
timestamp 1669390400
transform -1 0 70448 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__CLK
timestamp 1669390400
transform 1 0 53648 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__CLK
timestamp 1669390400
transform -1 0 54208 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__CLK
timestamp 1669390400
transform 1 0 52640 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__CLK
timestamp 1669390400
transform 1 0 56560 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__CLK
timestamp 1669390400
transform 1 0 54880 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__CLK
timestamp 1669390400
transform -1 0 81424 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__CLK
timestamp 1669390400
transform 1 0 76496 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__CLK
timestamp 1669390400
transform 1 0 87584 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__CLK
timestamp 1669390400
transform -1 0 88816 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__CLK
timestamp 1669390400
transform 1 0 82208 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__CLK
timestamp 1669390400
transform 1 0 88928 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__CLK
timestamp 1669390400
transform 1 0 67536 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__CLK
timestamp 1669390400
transform 1 0 79856 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__CLK
timestamp 1669390400
transform -1 0 53984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__CLK
timestamp 1669390400
transform 1 0 68320 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__CLK
timestamp 1669390400
transform 1 0 53760 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__CLK
timestamp 1669390400
transform 1 0 57344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__CLK
timestamp 1669390400
transform 1 0 53312 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1922__CLK
timestamp 1669390400
transform 1 0 58576 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__CLK
timestamp 1669390400
transform 1 0 76160 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__CLK
timestamp 1669390400
transform 1 0 57792 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__CLK
timestamp 1669390400
transform 1 0 76048 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1669390400
transform 1 0 83216 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1669390400
transform 1 0 62048 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1669390400
transform 1 0 88256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1669390400
transform 1 0 63168 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1669390400
transform 1 0 86576 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_clk_I
timestamp 1669390400
transform 1 0 58128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_clk_I
timestamp 1669390400
transform -1 0 64848 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_clk_I
timestamp 1669390400
transform 1 0 61376 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_clk_I
timestamp 1669390400
transform 1 0 60592 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_clk_I
timestamp 1669390400
transform 1 0 64960 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_clk_I
timestamp 1669390400
transform 1 0 60592 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_clk_I
timestamp 1669390400
transform 1 0 55776 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_clk_I
timestamp 1669390400
transform 1 0 59248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_clk_I
timestamp 1669390400
transform 1 0 57680 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_clk_I
timestamp 1669390400
transform 1 0 56896 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_clk_I
timestamp 1669390400
transform 1 0 64288 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_clk_I
timestamp 1669390400
transform 1 0 62048 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_clk_I
timestamp 1669390400
transform -1 0 66416 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_clk_I
timestamp 1669390400
transform 1 0 69664 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_clk_I
timestamp 1669390400
transform 1 0 62944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_clk_I
timestamp 1669390400
transform 1 0 69216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_clk_I
timestamp 1669390400
transform 1 0 82992 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_clk_I
timestamp 1669390400
transform 1 0 84448 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_clk_I
timestamp 1669390400
transform 1 0 84112 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_clk_I
timestamp 1669390400
transform 1 0 83440 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_clk_I
timestamp 1669390400
transform 1 0 90944 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_clk_I
timestamp 1669390400
transform 1 0 93072 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_clk_I
timestamp 1669390400
transform -1 0 95200 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_clk_I
timestamp 1669390400
transform 1 0 90608 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_24_clk_I
timestamp 1669390400
transform 1 0 90832 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_clk_I
timestamp 1669390400
transform 1 0 95536 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_clk_I
timestamp 1669390400
transform 1 0 91840 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_clk_I
timestamp 1669390400
transform 1 0 90608 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_28_clk_I
timestamp 1669390400
transform 1 0 96880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_clk_I
timestamp 1669390400
transform 1 0 88480 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_clk_I
timestamp 1669390400
transform -1 0 87584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_clk_I
timestamp 1669390400
transform 1 0 93744 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_clk_I
timestamp 1669390400
transform -1 0 97328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_clk_I
timestamp 1669390400
transform 1 0 97888 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_clk_I
timestamp 1669390400
transform 1 0 95872 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_clk_I
timestamp 1669390400
transform 1 0 97104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_clk_I
timestamp 1669390400
transform 1 0 97104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_clk_I
timestamp 1669390400
transform 1 0 98000 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_39_clk_I
timestamp 1669390400
transform 1 0 88480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_40_clk_I
timestamp 1669390400
transform -1 0 87024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_41_clk_I
timestamp 1669390400
transform 1 0 81200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_42_clk_I
timestamp 1669390400
transform 1 0 84672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_43_clk_I
timestamp 1669390400
transform 1 0 83776 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_44_clk_I
timestamp 1669390400
transform 1 0 69216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_45_clk_I
timestamp 1669390400
transform 1 0 61824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_46_clk_I
timestamp 1669390400
transform 1 0 68544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_47_clk_I
timestamp 1669390400
transform 1 0 66640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_48_clk_I
timestamp 1669390400
transform 1 0 61712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_50_clk_I
timestamp 1669390400
transform -1 0 61488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_51_clk_I
timestamp 1669390400
transform 1 0 56000 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_52_clk_I
timestamp 1669390400
transform 1 0 59920 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 1904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 1904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 1904 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform 1 0 1680 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 6272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 18704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 31136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 44352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform -1 0 56112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 67872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform -1 0 80864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform -1 0 93296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform -1 0 95872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1669390400
transform 1 0 8288 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1669390400
transform 1 0 21280 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1669390400
transform 1 0 33040 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1669390400
transform 1 0 46592 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform 1 0 58352 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1669390400
transform 1 0 70448 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1669390400
transform 1 0 82880 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1669390400
transform 1 0 93072 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41
timestamp 1669390400
transform 1 0 5936 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6272 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7168 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68
timestamp 1669390400
transform 1 0 8960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_142 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_150
timestamp 1669390400
transform 1 0 18144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_152
timestamp 1669390400
transform 1 0 18368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_155
timestamp 1669390400
transform 1 0 18704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_163
timestamp 1669390400
transform 1 0 19600 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171
timestamp 1669390400
transform 1 0 20496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_263
timestamp 1669390400
transform 1 0 30800 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_266
timestamp 1669390400
transform 1 0 31136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_274
timestamp 1669390400
transform 1 0 32032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_278
timestamp 1669390400
transform 1 0 32480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_368
timestamp 1669390400
transform 1 0 42560 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_376
timestamp 1669390400
transform 1 0 43456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_380
timestamp 1669390400
transform 1 0 43904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_394
timestamp 1669390400
transform 1 0 45472 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_410
timestamp 1669390400
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1669390400
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_473
timestamp 1669390400
transform 1 0 54320 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_481
timestamp 1669390400
transform 1 0 55216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_485
timestamp 1669390400
transform 1 0 55664 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_499
timestamp 1669390400
transform 1 0 57232 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_515
timestamp 1669390400
transform 1 0 59024 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_523
timestamp 1669390400
transform 1 0 59920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_578
timestamp 1669390400
transform 1 0 66080 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_586
timestamp 1669390400
transform 1 0 66976 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_590
timestamp 1669390400
transform 1 0 67424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_594
timestamp 1669390400
transform 1 0 67872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_607
timestamp 1669390400
transform 1 0 69328 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_623
timestamp 1669390400
transform 1 0 71120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_627
timestamp 1669390400
transform 1 0 71568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1669390400
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1669390400
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_699
timestamp 1669390400
transform 1 0 79632 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_702
timestamp 1669390400
transform 1 0 79968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_706
timestamp 1669390400
transform 1 0 80416 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_710
timestamp 1669390400
transform 1 0 80864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_718
timestamp 1669390400
transform 1 0 81760 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_734
timestamp 1669390400
transform 1 0 83552 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_737
timestamp 1669390400
transform 1 0 83888 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_769
timestamp 1669390400
transform 1 0 87472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_772
timestamp 1669390400
transform 1 0 87808 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_804
timestamp 1669390400
transform 1 0 91392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_807
timestamp 1669390400
transform 1 0 91728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_815
timestamp 1669390400
transform 1 0 92624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_821
timestamp 1669390400
transform 1 0 93296 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_829
timestamp 1669390400
transform 1 0 94192 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_837
timestamp 1669390400
transform 1 0 95088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1669390400
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_842
timestamp 1669390400
transform 1 0 95648 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_858
timestamp 1669390400
transform 1 0 97440 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1669390400
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1669390400
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_421
timestamp 1669390400
transform 1 0 48496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_492
timestamp 1669390400
transform 1 0 56448 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_563
timestamp 1669390400
transform 1 0 64400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1669390400
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_634
timestamp 1669390400
transform 1 0 72352 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1669390400
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_705
timestamp 1669390400
transform 1 0 80304 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1669390400
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_712
timestamp 1669390400
transform 1 0 81088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_776
timestamp 1669390400
transform 1 0 88256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_780
timestamp 1669390400
transform 1 0 88704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_783
timestamp 1669390400
transform 1 0 89040 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_847
timestamp 1669390400
transform 1 0 96208 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1669390400
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_854
timestamp 1669390400
transform 1 0 96992 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_862
timestamp 1669390400
transform 1 0 97888 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1669390400
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_456
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_527
timestamp 1669390400
transform 1 0 60368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1669390400
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_598
timestamp 1669390400
transform 1 0 68320 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1669390400
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_669
timestamp 1669390400
transform 1 0 76272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1669390400
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_740
timestamp 1669390400
transform 1 0 84224 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1669390400
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_747
timestamp 1669390400
transform 1 0 85008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_811
timestamp 1669390400
transform 1 0 92176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_815
timestamp 1669390400
transform 1 0 92624 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_818
timestamp 1669390400
transform 1 0 92960 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_850
timestamp 1669390400
transform 1 0 96544 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1669390400
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_705
timestamp 1669390400
transform 1 0 80304 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_709
timestamp 1669390400
transform 1 0 80752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_712
timestamp 1669390400
transform 1 0 81088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_776
timestamp 1669390400
transform 1 0 88256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_780
timestamp 1669390400
transform 1 0 88704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_783
timestamp 1669390400
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_847
timestamp 1669390400
transform 1 0 96208 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1669390400
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_854
timestamp 1669390400
transform 1 0 96992 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_862
timestamp 1669390400
transform 1 0 97888 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1669390400
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1669390400
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1669390400
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1669390400
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1669390400
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1669390400
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1669390400
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1669390400
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_818
timestamp 1669390400
transform 1 0 92960 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_850
timestamp 1669390400
transform 1 0 96544 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1669390400
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1669390400
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1669390400
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1669390400
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1669390400
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1669390400
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1669390400
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1669390400
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1669390400
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_854
timestamp 1669390400
transform 1 0 96992 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_862
timestamp 1669390400
transform 1 0 97888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1669390400
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1669390400
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1669390400
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1669390400
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1669390400
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1669390400
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1669390400
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1669390400
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_818
timestamp 1669390400
transform 1 0 92960 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_850
timestamp 1669390400
transform 1 0 96544 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1669390400
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1669390400
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1669390400
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1669390400
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1669390400
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1669390400
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1669390400
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1669390400
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1669390400
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_854
timestamp 1669390400
transform 1 0 96992 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_862
timestamp 1669390400
transform 1 0 97888 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1669390400
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1669390400
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1669390400
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1669390400
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1669390400
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1669390400
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_818
timestamp 1669390400
transform 1 0 92960 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_850
timestamp 1669390400
transform 1 0 96544 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1669390400
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1669390400
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1669390400
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1669390400
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1669390400
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1669390400
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1669390400
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1669390400
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_854
timestamp 1669390400
transform 1 0 96992 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_862
timestamp 1669390400
transform 1 0 97888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1669390400
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1669390400
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1669390400
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1669390400
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1669390400
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1669390400
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_818
timestamp 1669390400
transform 1 0 92960 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_850
timestamp 1669390400
transform 1 0 96544 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_5
timestamp 1669390400
transform 1 0 1904 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_69
timestamp 1669390400
transform 1 0 9072 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1669390400
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1669390400
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1669390400
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1669390400
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1669390400
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1669390400
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1669390400
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1669390400
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_854
timestamp 1669390400
transform 1 0 96992 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_862
timestamp 1669390400
transform 1 0 97888 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_9
timestamp 1669390400
transform 1 0 2352 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_25
timestamp 1669390400
transform 1 0 4144 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_33
timestamp 1669390400
transform 1 0 5040 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1669390400
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1669390400
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1669390400
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1669390400
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1669390400
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1669390400
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1669390400
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_818
timestamp 1669390400
transform 1 0 92960 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_850
timestamp 1669390400
transform 1 0 96544 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1669390400
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1669390400
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1669390400
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1669390400
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1669390400
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1669390400
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1669390400
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1669390400
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1669390400
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_854
timestamp 1669390400
transform 1 0 96992 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_862
timestamp 1669390400
transform 1 0 97888 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1669390400
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1669390400
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1669390400
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1669390400
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1669390400
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1669390400
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1669390400
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1669390400
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_818
timestamp 1669390400
transform 1 0 92960 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_850
timestamp 1669390400
transform 1 0 96544 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1669390400
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1669390400
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1669390400
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1669390400
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1669390400
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1669390400
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1669390400
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1669390400
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_854
timestamp 1669390400
transform 1 0 96992 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_862
timestamp 1669390400
transform 1 0 97888 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1669390400
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1669390400
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1669390400
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1669390400
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1669390400
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1669390400
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1669390400
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_818
timestamp 1669390400
transform 1 0 92960 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_850
timestamp 1669390400
transform 1 0 96544 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1669390400
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1669390400
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1669390400
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1669390400
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1669390400
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1669390400
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1669390400
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1669390400
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_854
timestamp 1669390400
transform 1 0 96992 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_862
timestamp 1669390400
transform 1 0 97888 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1669390400
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1669390400
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1669390400
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1669390400
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1669390400
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1669390400
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1669390400
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1669390400
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_818
timestamp 1669390400
transform 1 0 92960 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_850
timestamp 1669390400
transform 1 0 96544 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1669390400
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1669390400
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1669390400
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1669390400
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1669390400
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1669390400
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1669390400
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1669390400
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_854
timestamp 1669390400
transform 1 0 96992 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_862
timestamp 1669390400
transform 1 0 97888 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1669390400
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1669390400
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1669390400
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1669390400
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1669390400
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1669390400
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1669390400
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_818
timestamp 1669390400
transform 1 0 92960 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_850
timestamp 1669390400
transform 1 0 96544 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1669390400
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1669390400
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1669390400
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1669390400
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1669390400
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1669390400
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1669390400
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1669390400
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_854
timestamp 1669390400
transform 1 0 96992 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_862
timestamp 1669390400
transform 1 0 97888 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1669390400
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1669390400
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1669390400
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1669390400
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1669390400
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1669390400
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1669390400
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_818
timestamp 1669390400
transform 1 0 92960 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_850
timestamp 1669390400
transform 1 0 96544 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1669390400
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1669390400
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1669390400
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1669390400
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1669390400
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1669390400
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1669390400
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1669390400
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_854
timestamp 1669390400
transform 1 0 96992 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_862
timestamp 1669390400
transform 1 0 97888 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1669390400
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1669390400
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1669390400
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1669390400
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1669390400
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1669390400
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_818
timestamp 1669390400
transform 1 0 92960 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_850
timestamp 1669390400
transform 1 0 96544 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1669390400
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1669390400
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1669390400
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1669390400
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1669390400
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1669390400
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1669390400
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1669390400
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_854
timestamp 1669390400
transform 1 0 96992 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_862
timestamp 1669390400
transform 1 0 97888 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1669390400
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1669390400
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1669390400
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1669390400
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1669390400
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1669390400
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1669390400
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_818
timestamp 1669390400
transform 1 0 92960 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_850
timestamp 1669390400
transform 1 0 96544 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1669390400
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1669390400
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1669390400
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1669390400
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1669390400
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1669390400
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1669390400
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1669390400
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_854
timestamp 1669390400
transform 1 0 96992 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_862
timestamp 1669390400
transform 1 0 97888 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1669390400
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1669390400
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1669390400
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1669390400
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1669390400
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1669390400
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_818
timestamp 1669390400
transform 1 0 92960 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_840
timestamp 1669390400
transform 1 0 95424 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_844
timestamp 1669390400
transform 1 0 95872 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_860
timestamp 1669390400
transform 1 0 97664 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_864
timestamp 1669390400
transform 1 0 98112 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1669390400
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1669390400
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1669390400
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1669390400
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1669390400
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1669390400
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1669390400
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1669390400
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_854
timestamp 1669390400
transform 1 0 96992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_862
timestamp 1669390400
transform 1 0 97888 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1669390400
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1669390400
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1669390400
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1669390400
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1669390400
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1669390400
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1669390400
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_818
timestamp 1669390400
transform 1 0 92960 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_850
timestamp 1669390400
transform 1 0 96544 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1669390400
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1669390400
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1669390400
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1669390400
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1669390400
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1669390400
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1669390400
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1669390400
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_854
timestamp 1669390400
transform 1 0 96992 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_862
timestamp 1669390400
transform 1 0 97888 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1669390400
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1669390400
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1669390400
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1669390400
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1669390400
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1669390400
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_818
timestamp 1669390400
transform 1 0 92960 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_850
timestamp 1669390400
transform 1 0 96544 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1669390400
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1669390400
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_712
timestamp 1669390400
transform 1 0 81088 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_728
timestamp 1669390400
transform 1 0 82880 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_732
timestamp 1669390400
transform 1 0 83328 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_736
timestamp 1669390400
transform 1 0 83776 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_753
timestamp 1669390400
transform 1 0 85680 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_769
timestamp 1669390400
transform 1 0 87472 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_777
timestamp 1669390400
transform 1 0 88368 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1669390400
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1669390400
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1669390400
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_854
timestamp 1669390400
transform 1 0 96992 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_862
timestamp 1669390400
transform 1 0 97888 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1669390400
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1669390400
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1669390400
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1669390400
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1669390400
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1669390400
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1669390400
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_818
timestamp 1669390400
transform 1 0 92960 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_850
timestamp 1669390400
transform 1 0 96544 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_602
timestamp 1669390400
transform 1 0 68768 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_606
timestamp 1669390400
transform 1 0 69216 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_614
timestamp 1669390400
transform 1 0 70112 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_616
timestamp 1669390400
transform 1 0 70336 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_619
timestamp 1669390400
transform 1 0 70672 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_635
timestamp 1669390400
transform 1 0 72464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1669390400
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1669390400
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_712
timestamp 1669390400
transform 1 0 81088 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_728
timestamp 1669390400
transform 1 0 82880 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_758
timestamp 1669390400
transform 1 0 86240 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_774
timestamp 1669390400
transform 1 0 88032 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_778
timestamp 1669390400
transform 1 0 88480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1669390400
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1669390400
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1669390400
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1669390400
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_854
timestamp 1669390400
transform 1 0 96992 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_862
timestamp 1669390400
transform 1 0 97888 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_479
timestamp 1669390400
transform 1 0 54992 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_489
timestamp 1669390400
transform 1 0 56112 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_493
timestamp 1669390400
transform 1 0 56560 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_495
timestamp 1669390400
transform 1 0 56784 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_498
timestamp 1669390400
transform 1 0 57120 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_502
timestamp 1669390400
transform 1 0 57568 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_506
timestamp 1669390400
transform 1 0 58016 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_522
timestamp 1669390400
transform 1 0 59808 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_530
timestamp 1669390400
transform 1 0 60704 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_537
timestamp 1669390400
transform 1 0 61488 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_569
timestamp 1669390400
transform 1 0 65072 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_577
timestamp 1669390400
transform 1 0 65968 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_581
timestamp 1669390400
transform 1 0 66416 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_588
timestamp 1669390400
transform 1 0 67200 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_590
timestamp 1669390400
transform 1 0 67424 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_597
timestamp 1669390400
transform 1 0 68208 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_599
timestamp 1669390400
transform 1 0 68432 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_612
timestamp 1669390400
transform 1 0 69888 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_614
timestamp 1669390400
transform 1 0 70112 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_617
timestamp 1669390400
transform 1 0 70448 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_648
timestamp 1669390400
transform 1 0 73920 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_664
timestamp 1669390400
transform 1 0 75712 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_668
timestamp 1669390400
transform 1 0 76160 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_671
timestamp 1669390400
transform 1 0 76496 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1669390400
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_708
timestamp 1669390400
transform 1 0 80640 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_724
timestamp 1669390400
transform 1 0 82432 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_732
timestamp 1669390400
transform 1 0 83328 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_734
timestamp 1669390400
transform 1 0 83552 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_741
timestamp 1669390400
transform 1 0 84336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_747
timestamp 1669390400
transform 1 0 85008 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_765
timestamp 1669390400
transform 1 0 87024 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_781
timestamp 1669390400
transform 1 0 88816 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_783
timestamp 1669390400
transform 1 0 89040 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_786
timestamp 1669390400
transform 1 0 89376 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_794
timestamp 1669390400
transform 1 0 90272 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_810
timestamp 1669390400
transform 1 0 92064 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_814
timestamp 1669390400
transform 1 0 92512 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_818
timestamp 1669390400
transform 1 0 92960 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_850
timestamp 1669390400
transform 1 0 96544 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_460
timestamp 1669390400
transform 1 0 52864 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_464
timestamp 1669390400
transform 1 0 53312 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_466
timestamp 1669390400
transform 1 0 53536 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_469
timestamp 1669390400
transform 1 0 53872 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_479
timestamp 1669390400
transform 1 0 54992 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_506
timestamp 1669390400
transform 1 0 58016 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_510
timestamp 1669390400
transform 1 0 58464 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_518
timestamp 1669390400
transform 1 0 59360 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_520
timestamp 1669390400
transform 1 0 59584 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_523
timestamp 1669390400
transform 1 0 59920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_527
timestamp 1669390400
transform 1 0 60368 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_531
timestamp 1669390400
transform 1 0 60816 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_535
timestamp 1669390400
transform 1 0 61264 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_552
timestamp 1669390400
transform 1 0 63168 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_556
timestamp 1669390400
transform 1 0 63616 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_564
timestamp 1669390400
transform 1 0 64512 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_572
timestamp 1669390400
transform 1 0 65408 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_602
timestamp 1669390400
transform 1 0 68768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_619
timestamp 1669390400
transform 1 0 70672 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_623
timestamp 1669390400
transform 1 0 71120 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_627
timestamp 1669390400
transform 1 0 71568 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_629
timestamp 1669390400
transform 1 0 71792 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_644
timestamp 1669390400
transform 1 0 73472 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_648
timestamp 1669390400
transform 1 0 73920 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_652
timestamp 1669390400
transform 1 0 74368 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_656
timestamp 1669390400
transform 1 0 74816 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_659
timestamp 1669390400
transform 1 0 75152 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_663
timestamp 1669390400
transform 1 0 75600 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_669
timestamp 1669390400
transform 1 0 76272 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_686
timestamp 1669390400
transform 1 0 78176 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_702
timestamp 1669390400
transform 1 0 79968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_706
timestamp 1669390400
transform 1 0 80416 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1669390400
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_712
timestamp 1669390400
transform 1 0 81088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_719
timestamp 1669390400
transform 1 0 81872 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_750
timestamp 1669390400
transform 1 0 85344 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_754
timestamp 1669390400
transform 1 0 85792 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_758
timestamp 1669390400
transform 1 0 86240 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_775
timestamp 1669390400
transform 1 0 88144 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_779
timestamp 1669390400
transform 1 0 88592 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_783
timestamp 1669390400
transform 1 0 89040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_786
timestamp 1669390400
transform 1 0 89376 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_803
timestamp 1669390400
transform 1 0 91280 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_807
timestamp 1669390400
transform 1 0 91728 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_823
timestamp 1669390400
transform 1 0 93520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_827
timestamp 1669390400
transform 1 0 93968 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_830
timestamp 1669390400
transform 1 0 94304 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_834
timestamp 1669390400
transform 1 0 94752 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1669390400
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_854
timestamp 1669390400
transform 1 0 96992 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_862
timestamp 1669390400
transform 1 0 97888 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_424
timestamp 1669390400
transform 1 0 48832 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_440
timestamp 1669390400
transform 1 0 50624 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_444
timestamp 1669390400
transform 1 0 51072 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_451
timestamp 1669390400
transform 1 0 51856 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_459
timestamp 1669390400
transform 1 0 52752 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_466
timestamp 1669390400
transform 1 0 53536 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_470
timestamp 1669390400
transform 1 0 53984 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_472
timestamp 1669390400
transform 1 0 54208 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_502
timestamp 1669390400
transform 1 0 57568 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_519
timestamp 1669390400
transform 1 0 59472 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_523
timestamp 1669390400
transform 1 0 59920 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_537
timestamp 1669390400
transform 1 0 61488 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_570
timestamp 1669390400
transform 1 0 65184 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_572
timestamp 1669390400
transform 1 0 65408 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_638
timestamp 1669390400
transform 1 0 72800 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_642
timestamp 1669390400
transform 1 0 73248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_646
timestamp 1669390400
transform 1 0 73696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_658
timestamp 1669390400
transform 1 0 75040 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_662
timestamp 1669390400
transform 1 0 75488 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_671
timestamp 1669390400
transform 1 0 76496 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1669390400
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_683
timestamp 1669390400
transform 1 0 77840 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_714
timestamp 1669390400
transform 1 0 81312 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_731
timestamp 1669390400
transform 1 0 83216 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_739
timestamp 1669390400
transform 1 0 84112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_743
timestamp 1669390400
transform 1 0 84560 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_747
timestamp 1669390400
transform 1 0 85008 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_751
timestamp 1669390400
transform 1 0 85456 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_781
timestamp 1669390400
transform 1 0 88816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_785
timestamp 1669390400
transform 1 0 89264 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1669390400
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_818
timestamp 1669390400
transform 1 0 92960 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_826
timestamp 1669390400
transform 1 0 93856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_830
timestamp 1669390400
transform 1 0 94304 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_860
timestamp 1669390400
transform 1 0 97664 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_864
timestamp 1669390400
transform 1 0 98112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_436
timestamp 1669390400
transform 1 0 50176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_440
timestamp 1669390400
transform 1 0 50624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_448
timestamp 1669390400
transform 1 0 51520 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_465
timestamp 1669390400
transform 1 0 53424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_529
timestamp 1669390400
transform 1 0 60592 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_560
timestamp 1669390400
transform 1 0 64064 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_566
timestamp 1669390400
transform 1 0 64736 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_577
timestamp 1669390400
transform 1 0 65968 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_581
timestamp 1669390400
transform 1 0 66416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_635
timestamp 1669390400
transform 1 0 72464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_657
timestamp 1669390400
transform 1 0 74928 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_661
timestamp 1669390400
transform 1 0 75376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_694
timestamp 1669390400
transform 1 0 79072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_696
timestamp 1669390400
transform 1 0 79296 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_703
timestamp 1669390400
transform 1 0 80080 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_707
timestamp 1669390400
transform 1 0 80528 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1669390400
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_712
timestamp 1669390400
transform 1 0 81088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_763
timestamp 1669390400
transform 1 0 86800 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1669390400
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_783
timestamp 1669390400
transform 1 0 89040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_813
timestamp 1669390400
transform 1 0 92400 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_821
timestamp 1669390400
transform 1 0 93296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_823
timestamp 1669390400
transform 1 0 93520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_826
timestamp 1669390400
transform 1 0 93856 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_834
timestamp 1669390400
transform 1 0 94752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1669390400
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_854
timestamp 1669390400
transform 1 0 96992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_857
timestamp 1669390400
transform 1 0 97328 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_865
timestamp 1669390400
transform 1 0 98224 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_424
timestamp 1669390400
transform 1 0 48832 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_428
timestamp 1669390400
transform 1 0 49280 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_430
timestamp 1669390400
transform 1 0 49504 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_466
timestamp 1669390400
transform 1 0 53536 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_470
timestamp 1669390400
transform 1 0 53984 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_478
timestamp 1669390400
transform 1 0 54880 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_480
timestamp 1669390400
transform 1 0 55104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_564
timestamp 1669390400
transform 1 0 64512 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_581
timestamp 1669390400
transform 1 0 66416 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_585
timestamp 1669390400
transform 1 0 66864 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_608
timestamp 1669390400
transform 1 0 69440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_612
timestamp 1669390400
transform 1 0 69888 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_616
timestamp 1669390400
transform 1 0 70336 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_618
timestamp 1669390400
transform 1 0 70560 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_625
timestamp 1669390400
transform 1 0 71344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_642
timestamp 1669390400
transform 1 0 73248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1669390400
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_679
timestamp 1669390400
transform 1 0 77392 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_687
timestamp 1669390400
transform 1 0 78288 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_689
timestamp 1669390400
transform 1 0 78512 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_719
timestamp 1669390400
transform 1 0 81872 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_736
timestamp 1669390400
transform 1 0 83776 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1669390400
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_747
timestamp 1669390400
transform 1 0 85008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_777
timestamp 1669390400
transform 1 0 88368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_781
timestamp 1669390400
transform 1 0 88816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_791
timestamp 1669390400
transform 1 0 89936 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_795
timestamp 1669390400
transform 1 0 90384 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_812
timestamp 1669390400
transform 1 0 92288 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_818
timestamp 1669390400
transform 1 0 92960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_826
timestamp 1669390400
transform 1 0 93856 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_828
timestamp 1669390400
transform 1 0 94080 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_858
timestamp 1669390400
transform 1 0 97440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_432
timestamp 1669390400
transform 1 0 49728 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_462
timestamp 1669390400
transform 1 0 53088 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_479
timestamp 1669390400
transform 1 0 54992 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_483
timestamp 1669390400
transform 1 0 55440 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_491
timestamp 1669390400
transform 1 0 56336 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_493
timestamp 1669390400
transform 1 0 56560 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_518
timestamp 1669390400
transform 1 0 59360 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_522
timestamp 1669390400
transform 1 0 59808 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_524
timestamp 1669390400
transform 1 0 60032 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_531
timestamp 1669390400
transform 1 0 60816 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_535
timestamp 1669390400
transform 1 0 61264 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_554
timestamp 1669390400
transform 1 0 63392 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_558
timestamp 1669390400
transform 1 0 63840 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_562
timestamp 1669390400
transform 1 0 64288 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_566
timestamp 1669390400
transform 1 0 64736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_578
timestamp 1669390400
transform 1 0 66080 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_582
timestamp 1669390400
transform 1 0 66528 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_585
timestamp 1669390400
transform 1 0 66864 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_617
timestamp 1669390400
transform 1 0 70448 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_625
timestamp 1669390400
transform 1 0 71344 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_633
timestamp 1669390400
transform 1 0 72240 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_635
timestamp 1669390400
transform 1 0 72464 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_651
timestamp 1669390400
transform 1 0 74256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_668
timestamp 1669390400
transform 1 0 76160 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_676
timestamp 1669390400
transform 1 0 77056 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_680
timestamp 1669390400
transform 1 0 77504 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_696
timestamp 1669390400
transform 1 0 79296 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_704
timestamp 1669390400
transform 1 0 80192 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_708
timestamp 1669390400
transform 1 0 80640 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_712
timestamp 1669390400
transform 1 0 81088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_715
timestamp 1669390400
transform 1 0 81424 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_719
timestamp 1669390400
transform 1 0 81872 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_723
timestamp 1669390400
transform 1 0 82320 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_726
timestamp 1669390400
transform 1 0 82656 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_734
timestamp 1669390400
transform 1 0 83552 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_744
timestamp 1669390400
transform 1 0 84672 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_748
timestamp 1669390400
transform 1 0 85120 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_765
timestamp 1669390400
transform 1 0 87024 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_775
timestamp 1669390400
transform 1 0 88144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_777
timestamp 1669390400
transform 1 0 88368 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1669390400
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_783
timestamp 1669390400
transform 1 0 89040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_799
timestamp 1669390400
transform 1 0 90832 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1669390400
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_854
timestamp 1669390400
transform 1 0 96992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_857
timestamp 1669390400
transform 1 0 97328 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_865
timestamp 1669390400
transform 1 0 98224 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_424
timestamp 1669390400
transform 1 0 48832 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_440
timestamp 1669390400
transform 1 0 50624 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_457
timestamp 1669390400
transform 1 0 52528 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_466
timestamp 1669390400
transform 1 0 53536 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_470
timestamp 1669390400
transform 1 0 53984 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_474
timestamp 1669390400
transform 1 0 54432 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_482
timestamp 1669390400
transform 1 0 55328 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_486
timestamp 1669390400
transform 1 0 55776 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_516
timestamp 1669390400
transform 1 0 59136 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_524
timestamp 1669390400
transform 1 0 60032 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_528
timestamp 1669390400
transform 1 0 60480 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_534
timestamp 1669390400
transform 1 0 61152 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_536
timestamp 1669390400
transform 1 0 61376 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_539
timestamp 1669390400
transform 1 0 61712 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_555
timestamp 1669390400
transform 1 0 63504 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_563
timestamp 1669390400
transform 1 0 64400 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_569
timestamp 1669390400
transform 1 0 65072 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_573
timestamp 1669390400
transform 1 0 65520 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_589
timestamp 1669390400
transform 1 0 67312 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_593
timestamp 1669390400
transform 1 0 67760 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_600
timestamp 1669390400
transform 1 0 68544 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1669390400
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_605
timestamp 1669390400
transform 1 0 69104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_621
timestamp 1669390400
transform 1 0 70896 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_625
timestamp 1669390400
transform 1 0 71344 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_629
timestamp 1669390400
transform 1 0 71792 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_637
timestamp 1669390400
transform 1 0 72688 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_641
timestamp 1669390400
transform 1 0 73136 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_644
timestamp 1669390400
transform 1 0 73472 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_654
timestamp 1669390400
transform 1 0 74592 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_664
timestamp 1669390400
transform 1 0 75712 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_672
timestamp 1669390400
transform 1 0 76608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_676
timestamp 1669390400
transform 1 0 77056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_679
timestamp 1669390400
transform 1 0 77392 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_683
timestamp 1669390400
transform 1 0 77840 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_715
timestamp 1669390400
transform 1 0 81424 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_723
timestamp 1669390400
transform 1 0 82320 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_726
timestamp 1669390400
transform 1 0 82656 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_742
timestamp 1669390400
transform 1 0 84448 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_744
timestamp 1669390400
transform 1 0 84672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_747
timestamp 1669390400
transform 1 0 85008 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_763
timestamp 1669390400
transform 1 0 86800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_767
timestamp 1669390400
transform 1 0 87248 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_783
timestamp 1669390400
transform 1 0 89040 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_785
timestamp 1669390400
transform 1 0 89264 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_815
timestamp 1669390400
transform 1 0 92624 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_818
timestamp 1669390400
transform 1 0 92960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_822
timestamp 1669390400
transform 1 0 93408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_826
timestamp 1669390400
transform 1 0 93856 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_834
timestamp 1669390400
transform 1 0 94752 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_851
timestamp 1669390400
transform 1 0 96656 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_855
timestamp 1669390400
transform 1 0 97104 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_863
timestamp 1669390400
transform 1 0 98000 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_865
timestamp 1669390400
transform 1 0 98224 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_5
timestamp 1669390400
transform 1 0 1904 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_69
timestamp 1669390400
transform 1 0 9072 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_458
timestamp 1669390400
transform 1 0 52640 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_462
timestamp 1669390400
transform 1 0 53088 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_478
timestamp 1669390400
transform 1 0 54880 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_486
timestamp 1669390400
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_516
timestamp 1669390400
transform 1 0 59136 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_520
timestamp 1669390400
transform 1 0 59584 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_524
timestamp 1669390400
transform 1 0 60032 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_540
timestamp 1669390400
transform 1 0 61824 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_548
timestamp 1669390400
transform 1 0 62720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1669390400
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_570
timestamp 1669390400
transform 1 0 65184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_573
timestamp 1669390400
transform 1 0 65520 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_577
timestamp 1669390400
transform 1 0 65968 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_581
timestamp 1669390400
transform 1 0 66416 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_611
timestamp 1669390400
transform 1 0 69776 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_615
timestamp 1669390400
transform 1 0 70224 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_631
timestamp 1669390400
transform 1 0 72016 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_641
timestamp 1669390400
transform 1 0 73136 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_649
timestamp 1669390400
transform 1 0 74032 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_652
timestamp 1669390400
transform 1 0 74368 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_656
timestamp 1669390400
transform 1 0 74816 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_673
timestamp 1669390400
transform 1 0 76720 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_677
timestamp 1669390400
transform 1 0 77168 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_681
timestamp 1669390400
transform 1 0 77616 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_685
timestamp 1669390400
transform 1 0 78064 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_701
timestamp 1669390400
transform 1 0 79856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_709
timestamp 1669390400
transform 1 0 80752 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_712
timestamp 1669390400
transform 1 0 81088 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_716
timestamp 1669390400
transform 1 0 81536 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_724
timestamp 1669390400
transform 1 0 82432 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_741
timestamp 1669390400
transform 1 0 84336 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_745
timestamp 1669390400
transform 1 0 84784 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_777
timestamp 1669390400
transform 1 0 88368 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_783
timestamp 1669390400
transform 1 0 89040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_813
timestamp 1669390400
transform 1 0 92400 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_821
timestamp 1669390400
transform 1 0 93296 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_827
timestamp 1669390400
transform 1 0 93968 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_831
timestamp 1669390400
transform 1 0 94416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_835
timestamp 1669390400
transform 1 0 94864 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_851
timestamp 1669390400
transform 1 0 96656 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_854
timestamp 1669390400
transform 1 0 96992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_857
timestamp 1669390400
transform 1 0 97328 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_865
timestamp 1669390400
transform 1 0 98224 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_9
timestamp 1669390400
transform 1 0 2352 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_25
timestamp 1669390400
transform 1 0 4144 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_33
timestamp 1669390400
transform 1 0 5040 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_408
timestamp 1669390400
transform 1 0 47040 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_416
timestamp 1669390400
transform 1 0 47936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_420
timestamp 1669390400
transform 1 0 48384 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_422
timestamp 1669390400
transform 1 0 48608 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_429
timestamp 1669390400
transform 1 0 49392 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_466
timestamp 1669390400
transform 1 0 53536 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_470
timestamp 1669390400
transform 1 0 53984 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_478
timestamp 1669390400
transform 1 0 54880 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_482
timestamp 1669390400
transform 1 0 55328 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_484
timestamp 1669390400
transform 1 0 55552 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_487
timestamp 1669390400
transform 1 0 55888 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_504
timestamp 1669390400
transform 1 0 57792 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_508
timestamp 1669390400
transform 1 0 58240 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_524
timestamp 1669390400
transform 1 0 60032 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_534
timestamp 1669390400
transform 1 0 61152 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_536
timestamp 1669390400
transform 1 0 61376 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_539
timestamp 1669390400
transform 1 0 61712 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_570
timestamp 1669390400
transform 1 0 65184 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_574
timestamp 1669390400
transform 1 0 65632 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_584
timestamp 1669390400
transform 1 0 66752 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_601
timestamp 1669390400
transform 1 0 68656 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_605
timestamp 1669390400
transform 1 0 69104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_608
timestamp 1669390400
transform 1 0 69440 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_612
timestamp 1669390400
transform 1 0 69888 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_644
timestamp 1669390400
transform 1 0 73472 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_652
timestamp 1669390400
transform 1 0 74368 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_669
timestamp 1669390400
transform 1 0 76272 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1669390400
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_676
timestamp 1669390400
transform 1 0 77056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_685
timestamp 1669390400
transform 1 0 78064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_691
timestamp 1669390400
transform 1 0 78736 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_695
timestamp 1669390400
transform 1 0 79184 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_711
timestamp 1669390400
transform 1 0 80976 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_742
timestamp 1669390400
transform 1 0 84448 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_744
timestamp 1669390400
transform 1 0 84672 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_747
timestamp 1669390400
transform 1 0 85008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_750
timestamp 1669390400
transform 1 0 85344 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_766
timestamp 1669390400
transform 1 0 87136 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_774
timestamp 1669390400
transform 1 0 88032 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_780
timestamp 1669390400
transform 1 0 88704 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_788
timestamp 1669390400
transform 1 0 89600 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_792
timestamp 1669390400
transform 1 0 90048 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_796
timestamp 1669390400
transform 1 0 90496 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_812
timestamp 1669390400
transform 1 0 92288 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_818
timestamp 1669390400
transform 1 0 92960 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_822
timestamp 1669390400
transform 1 0 93408 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_830
timestamp 1669390400
transform 1 0 94304 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_861
timestamp 1669390400
transform 1 0 97776 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_865
timestamp 1669390400
transform 1 0 98224 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_442
timestamp 1669390400
transform 1 0 50848 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_459
timestamp 1669390400
transform 1 0 52752 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_463
timestamp 1669390400
transform 1 0 53200 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_507
timestamp 1669390400
transform 1 0 58128 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_509
timestamp 1669390400
transform 1 0 58352 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_539
timestamp 1669390400
transform 1 0 61712 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_556
timestamp 1669390400
transform 1 0 63616 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_564
timestamp 1669390400
transform 1 0 64512 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_570
timestamp 1669390400
transform 1 0 65184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_600
timestamp 1669390400
transform 1 0 68544 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_623
timestamp 1669390400
transform 1 0 71120 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_627
timestamp 1669390400
transform 1 0 71568 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_631
timestamp 1669390400
transform 1 0 72016 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_641
timestamp 1669390400
transform 1 0 73136 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_649
timestamp 1669390400
transform 1 0 74032 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_651
timestamp 1669390400
transform 1 0 74256 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_658
timestamp 1669390400
transform 1 0 75040 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_689
timestamp 1669390400
transform 1 0 78512 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_706
timestamp 1669390400
transform 1 0 80416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_712
timestamp 1669390400
transform 1 0 81088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_715
timestamp 1669390400
transform 1 0 81424 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_752
timestamp 1669390400
transform 1 0 85568 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_756
timestamp 1669390400
transform 1 0 86016 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_772
timestamp 1669390400
transform 1 0 87808 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_776
timestamp 1669390400
transform 1 0 88256 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_780
timestamp 1669390400
transform 1 0 88704 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_783
timestamp 1669390400
transform 1 0 89040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_790
timestamp 1669390400
transform 1 0 89824 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_798
timestamp 1669390400
transform 1 0 90720 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_829
timestamp 1669390400
transform 1 0 94192 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_831
timestamp 1669390400
transform 1 0 94416 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_834
timestamp 1669390400
transform 1 0 94752 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_851
timestamp 1669390400
transform 1 0 96656 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_854
timestamp 1669390400
transform 1 0 96992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_857
timestamp 1669390400
transform 1 0 97328 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_861
timestamp 1669390400
transform 1 0 97776 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_865
timestamp 1669390400
transform 1 0 98224 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_424
timestamp 1669390400
transform 1 0 48832 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_432
timestamp 1669390400
transform 1 0 49728 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_436
timestamp 1669390400
transform 1 0 50176 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_438
timestamp 1669390400
transform 1 0 50400 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_441
timestamp 1669390400
transform 1 0 50736 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_449
timestamp 1669390400
transform 1 0 51632 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_457
timestamp 1669390400
transform 1 0 52528 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_467
timestamp 1669390400
transform 1 0 53648 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_475
timestamp 1669390400
transform 1 0 54544 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_479
timestamp 1669390400
transform 1 0 54992 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_481
timestamp 1669390400
transform 1 0 55216 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_488
timestamp 1669390400
transform 1 0 56000 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_504
timestamp 1669390400
transform 1 0 57792 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_512
timestamp 1669390400
transform 1 0 58688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_516
timestamp 1669390400
transform 1 0 59136 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_518
timestamp 1669390400
transform 1 0 59360 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_525
timestamp 1669390400
transform 1 0 60144 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_529
timestamp 1669390400
transform 1 0 60592 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1669390400
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_534
timestamp 1669390400
transform 1 0 61152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_537
timestamp 1669390400
transform 1 0 61488 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_541
timestamp 1669390400
transform 1 0 61936 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_593
timestamp 1669390400
transform 1 0 67760 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_595
timestamp 1669390400
transform 1 0 67984 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1669390400
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_605
timestamp 1669390400
transform 1 0 69104 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_617
timestamp 1669390400
transform 1 0 70448 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_621
timestamp 1669390400
transform 1 0 70896 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_658
timestamp 1669390400
transform 1 0 75040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_668
timestamp 1669390400
transform 1 0 76160 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_672
timestamp 1669390400
transform 1 0 76608 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_676
timestamp 1669390400
transform 1 0 77056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_679
timestamp 1669390400
transform 1 0 77392 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_685
timestamp 1669390400
transform 1 0 78064 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_716
timestamp 1669390400
transform 1 0 81536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_720
timestamp 1669390400
transform 1 0 81984 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_727
timestamp 1669390400
transform 1 0 82768 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_744
timestamp 1669390400
transform 1 0 84672 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_747
timestamp 1669390400
transform 1 0 85008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_750
timestamp 1669390400
transform 1 0 85344 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_766
timestamp 1669390400
transform 1 0 87136 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_770
timestamp 1669390400
transform 1 0 87584 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_801
timestamp 1669390400
transform 1 0 91056 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_809
timestamp 1669390400
transform 1 0 91952 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_813
timestamp 1669390400
transform 1 0 92400 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_815
timestamp 1669390400
transform 1 0 92624 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_818
timestamp 1669390400
transform 1 0 92960 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_820
timestamp 1669390400
transform 1 0 93184 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_823
timestamp 1669390400
transform 1 0 93520 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_831
timestamp 1669390400
transform 1 0 94416 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_833
timestamp 1669390400
transform 1 0 94640 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_863
timestamp 1669390400
transform 1 0 98000 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_865
timestamp 1669390400
transform 1 0 98224 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_66
timestamp 1669390400
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_421
timestamp 1669390400
transform 1 0 48496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1669390400
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_486
timestamp 1669390400
transform 1 0 55776 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_490
timestamp 1669390400
transform 1 0 56224 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_494
timestamp 1669390400
transform 1 0 56672 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_509
timestamp 1669390400
transform 1 0 58352 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_511
timestamp 1669390400
transform 1 0 58576 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_541
timestamp 1669390400
transform 1 0 61936 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_545
timestamp 1669390400
transform 1 0 62384 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_547
timestamp 1669390400
transform 1 0 62608 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_550
timestamp 1669390400
transform 1 0 62944 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1669390400
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_570
timestamp 1669390400
transform 1 0 65184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_573
timestamp 1669390400
transform 1 0 65520 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_581
timestamp 1669390400
transform 1 0 66416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_585
timestamp 1669390400
transform 1 0 66864 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_587
timestamp 1669390400
transform 1 0 67088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_617
timestamp 1669390400
transform 1 0 70448 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_621
timestamp 1669390400
transform 1 0 70896 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_631
timestamp 1669390400
transform 1 0 72016 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_635
timestamp 1669390400
transform 1 0 72464 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_641
timestamp 1669390400
transform 1 0 73136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_648
timestamp 1669390400
transform 1 0 73920 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_652
timestamp 1669390400
transform 1 0 74368 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_656
timestamp 1669390400
transform 1 0 74816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_708
timestamp 1669390400
transform 1 0 80640 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_712
timestamp 1669390400
transform 1 0 81088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_715
timestamp 1669390400
transform 1 0 81424 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_723
timestamp 1669390400
transform 1 0 82320 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_725
timestamp 1669390400
transform 1 0 82544 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_728
timestamp 1669390400
transform 1 0 82880 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_780
timestamp 1669390400
transform 1 0 88704 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_783
timestamp 1669390400
transform 1 0 89040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_790
timestamp 1669390400
transform 1 0 89824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_844
timestamp 1669390400
transform 1 0 95872 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_848
timestamp 1669390400
transform 1 0 96320 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_854
timestamp 1669390400
transform 1 0 96992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_861
timestamp 1669390400
transform 1 0 97776 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_865
timestamp 1669390400
transform 1 0 98224 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_424
timestamp 1669390400
transform 1 0 48832 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_428
timestamp 1669390400
transform 1 0 49280 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_435
timestamp 1669390400
transform 1 0 50064 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_443
timestamp 1669390400
transform 1 0 50960 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_466
timestamp 1669390400
transform 1 0 53536 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_470
timestamp 1669390400
transform 1 0 53984 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_474
timestamp 1669390400
transform 1 0 54432 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_478
timestamp 1669390400
transform 1 0 54880 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_482
timestamp 1669390400
transform 1 0 55328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_490
timestamp 1669390400
transform 1 0 56224 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_494
timestamp 1669390400
transform 1 0 56672 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_498
timestamp 1669390400
transform 1 0 57120 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_500
timestamp 1669390400
transform 1 0 57344 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_507
timestamp 1669390400
transform 1 0 58128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_524
timestamp 1669390400
transform 1 0 60032 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_528
timestamp 1669390400
transform 1 0 60480 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_534
timestamp 1669390400
transform 1 0 61152 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_571
timestamp 1669390400
transform 1 0 65296 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_575
timestamp 1669390400
transform 1 0 65744 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_579
timestamp 1669390400
transform 1 0 66192 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_587
timestamp 1669390400
transform 1 0 67088 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_594
timestamp 1669390400
transform 1 0 67872 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_598
timestamp 1669390400
transform 1 0 68320 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1669390400
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_605
timestamp 1669390400
transform 1 0 69104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_614
timestamp 1669390400
transform 1 0 70112 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_618
timestamp 1669390400
transform 1 0 70560 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_622
timestamp 1669390400
transform 1 0 71008 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_626
timestamp 1669390400
transform 1 0 71456 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_635
timestamp 1669390400
transform 1 0 72464 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_639
timestamp 1669390400
transform 1 0 72912 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_641
timestamp 1669390400
transform 1 0 73136 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_657
timestamp 1669390400
transform 1 0 74928 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_667
timestamp 1669390400
transform 1 0 76048 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_671
timestamp 1669390400
transform 1 0 76496 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1669390400
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_676
timestamp 1669390400
transform 1 0 77056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_683
timestamp 1669390400
transform 1 0 77840 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_691
timestamp 1669390400
transform 1 0 78736 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_698
timestamp 1669390400
transform 1 0 79520 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_714
timestamp 1669390400
transform 1 0 81312 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_717
timestamp 1669390400
transform 1 0 81648 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_734
timestamp 1669390400
transform 1 0 83552 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_738
timestamp 1669390400
transform 1 0 84000 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_742
timestamp 1669390400
transform 1 0 84448 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_744
timestamp 1669390400
transform 1 0 84672 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_747
timestamp 1669390400
transform 1 0 85008 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_757
timestamp 1669390400
transform 1 0 86128 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_790
timestamp 1669390400
transform 1 0 89824 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_807
timestamp 1669390400
transform 1 0 91728 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_815
timestamp 1669390400
transform 1 0 92624 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_818
timestamp 1669390400
transform 1 0 92960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_848
timestamp 1669390400
transform 1 0 96320 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_865
timestamp 1669390400
transform 1 0 98224 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_421
timestamp 1669390400
transform 1 0 48496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_458
timestamp 1669390400
transform 1 0 52640 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_475
timestamp 1669390400
transform 1 0 54544 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_479
timestamp 1669390400
transform 1 0 54992 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_550
timestamp 1669390400
transform 1 0 62944 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1669390400
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_570
timestamp 1669390400
transform 1 0 65184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_577
timestamp 1669390400
transform 1 0 65968 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_608
timestamp 1669390400
transform 1 0 69440 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_625
timestamp 1669390400
transform 1 0 71344 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_635
timestamp 1669390400
transform 1 0 72464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_641
timestamp 1669390400
transform 1 0 73136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_644
timestamp 1669390400
transform 1 0 73472 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_646
timestamp 1669390400
transform 1 0 73696 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_676
timestamp 1669390400
transform 1 0 77056 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_680
timestamp 1669390400
transform 1 0 77504 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_684
timestamp 1669390400
transform 1 0 77952 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_688
timestamp 1669390400
transform 1 0 78400 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_704
timestamp 1669390400
transform 1 0 80192 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_708
timestamp 1669390400
transform 1 0 80640 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_712
timestamp 1669390400
transform 1 0 81088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_742
timestamp 1669390400
transform 1 0 84448 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_773
timestamp 1669390400
transform 1 0 87920 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_777
timestamp 1669390400
transform 1 0 88368 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_783
timestamp 1669390400
transform 1 0 89040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_834
timestamp 1669390400
transform 1 0 94752 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_851
timestamp 1669390400
transform 1 0 96656 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_854
timestamp 1669390400
transform 1 0 96992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_861
timestamp 1669390400
transform 1 0 97776 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_865
timestamp 1669390400
transform 1 0 98224 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_424
timestamp 1669390400
transform 1 0 48832 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_428
timestamp 1669390400
transform 1 0 49280 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_430
timestamp 1669390400
transform 1 0 49504 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1669390400
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_466
timestamp 1669390400
transform 1 0 53536 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_468
timestamp 1669390400
transform 1 0 53760 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_498
timestamp 1669390400
transform 1 0 57120 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_529
timestamp 1669390400
transform 1 0 60592 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1669390400
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_534
timestamp 1669390400
transform 1 0 61152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_537
timestamp 1669390400
transform 1 0 61488 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_541
timestamp 1669390400
transform 1 0 61936 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_544
timestamp 1669390400
transform 1 0 62272 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_548
timestamp 1669390400
transform 1 0 62720 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_579
timestamp 1669390400
transform 1 0 66192 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_583
timestamp 1669390400
transform 1 0 66640 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_599
timestamp 1669390400
transform 1 0 68432 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1669390400
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_605
timestamp 1669390400
transform 1 0 69104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_656
timestamp 1669390400
transform 1 0 74816 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_666
timestamp 1669390400
transform 1 0 75936 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_670
timestamp 1669390400
transform 1 0 76384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_676
timestamp 1669390400
transform 1 0 77056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_692
timestamp 1669390400
transform 1 0 78848 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_696
timestamp 1669390400
transform 1 0 79296 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_712
timestamp 1669390400
transform 1 0 81088 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_722
timestamp 1669390400
transform 1 0 82208 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_738
timestamp 1669390400
transform 1 0 84000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_742
timestamp 1669390400
transform 1 0 84448 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_744
timestamp 1669390400
transform 1 0 84672 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_747
timestamp 1669390400
transform 1 0 85008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_750
timestamp 1669390400
transform 1 0 85344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_767
timestamp 1669390400
transform 1 0 87248 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_771
timestamp 1669390400
transform 1 0 87696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_775
timestamp 1669390400
transform 1 0 88144 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_778
timestamp 1669390400
transform 1 0 88480 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_782
timestamp 1669390400
transform 1 0 88928 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_799
timestamp 1669390400
transform 1 0 90832 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_807
timestamp 1669390400
transform 1 0 91728 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_811
timestamp 1669390400
transform 1 0 92176 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_815
timestamp 1669390400
transform 1 0 92624 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_818
timestamp 1669390400
transform 1 0 92960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_825
timestamp 1669390400
transform 1 0 93744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_829
timestamp 1669390400
transform 1 0 94192 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_832
timestamp 1669390400
transform 1 0 94528 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_863
timestamp 1669390400
transform 1 0 98000 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_865
timestamp 1669390400
transform 1 0 98224 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1669390400
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_405
timestamp 1669390400
transform 1 0 46704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_413
timestamp 1669390400
transform 1 0 47600 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_417
timestamp 1669390400
transform 1 0 48048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_445
timestamp 1669390400
transform 1 0 51184 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_462
timestamp 1669390400
transform 1 0 53088 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_466
timestamp 1669390400
transform 1 0 53536 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_470
timestamp 1669390400
transform 1 0 53984 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_474
timestamp 1669390400
transform 1 0 54432 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_484
timestamp 1669390400
transform 1 0 55552 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_515
timestamp 1669390400
transform 1 0 59024 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_519
timestamp 1669390400
transform 1 0 59472 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_527
timestamp 1669390400
transform 1 0 60368 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_543
timestamp 1669390400
transform 1 0 62160 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_551
timestamp 1669390400
transform 1 0 63056 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1669390400
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_570
timestamp 1669390400
transform 1 0 65184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_573
timestamp 1669390400
transform 1 0 65520 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_577
timestamp 1669390400
transform 1 0 65968 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_593
timestamp 1669390400
transform 1 0 67760 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_601
timestamp 1669390400
transform 1 0 68656 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_605
timestamp 1669390400
transform 1 0 69104 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_609
timestamp 1669390400
transform 1 0 69552 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_617
timestamp 1669390400
transform 1 0 70448 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_634
timestamp 1669390400
transform 1 0 72352 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1669390400
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_641
timestamp 1669390400
transform 1 0 73136 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_649
timestamp 1669390400
transform 1 0 74032 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_655
timestamp 1669390400
transform 1 0 74704 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_672
timestamp 1669390400
transform 1 0 76608 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_674
timestamp 1669390400
transform 1 0 76832 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_704
timestamp 1669390400
transform 1 0 80192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_708
timestamp 1669390400
transform 1 0 80640 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_712
timestamp 1669390400
transform 1 0 81088 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_746
timestamp 1669390400
transform 1 0 84896 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_778
timestamp 1669390400
transform 1 0 88480 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_780
timestamp 1669390400
transform 1 0 88704 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_783
timestamp 1669390400
transform 1 0 89040 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_787
timestamp 1669390400
transform 1 0 89488 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_790
timestamp 1669390400
transform 1 0 89824 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_794
timestamp 1669390400
transform 1 0 90272 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_798
timestamp 1669390400
transform 1 0 90720 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_800
timestamp 1669390400
transform 1 0 90944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_851
timestamp 1669390400
transform 1 0 96656 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_854
timestamp 1669390400
transform 1 0 96992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_857
timestamp 1669390400
transform 1 0 97328 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_865
timestamp 1669390400
transform 1 0 98224 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_385
timestamp 1669390400
transform 1 0 44464 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_453
timestamp 1669390400
transform 1 0 52080 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_457
timestamp 1669390400
transform 1 0 52528 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_479
timestamp 1669390400
transform 1 0 54992 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_509
timestamp 1669390400
transform 1 0 58352 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_513
timestamp 1669390400
transform 1 0 58800 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_519
timestamp 1669390400
transform 1 0 59472 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_527
timestamp 1669390400
transform 1 0 60368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1669390400
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_534
timestamp 1669390400
transform 1 0 61152 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_538
timestamp 1669390400
transform 1 0 61600 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_542
timestamp 1669390400
transform 1 0 62048 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_550
timestamp 1669390400
transform 1 0 62944 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1669390400
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_605
timestamp 1669390400
transform 1 0 69104 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_636
timestamp 1669390400
transform 1 0 72576 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_640
timestamp 1669390400
transform 1 0 73024 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1669390400
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_676
timestamp 1669390400
transform 1 0 77056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_692
timestamp 1669390400
transform 1 0 78848 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_744
timestamp 1669390400
transform 1 0 84672 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_747
timestamp 1669390400
transform 1 0 85008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_754
timestamp 1669390400
transform 1 0 85792 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_786
timestamp 1669390400
transform 1 0 89376 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_794
timestamp 1669390400
transform 1 0 90272 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_798
timestamp 1669390400
transform 1 0 90720 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_815
timestamp 1669390400
transform 1 0 92624 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_818
timestamp 1669390400
transform 1 0 92960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_821
timestamp 1669390400
transform 1 0 93296 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_825
timestamp 1669390400
transform 1 0 93744 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_829
timestamp 1669390400
transform 1 0 94192 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_833
timestamp 1669390400
transform 1 0 94640 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_863
timestamp 1669390400
transform 1 0 98000 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_865
timestamp 1669390400
transform 1 0 98224 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_432
timestamp 1669390400
transform 1 0 49728 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_462
timestamp 1669390400
transform 1 0 53088 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_466
timestamp 1669390400
transform 1 0 53536 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_482
timestamp 1669390400
transform 1 0 55328 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_486
timestamp 1669390400
transform 1 0 55776 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_488
timestamp 1669390400
transform 1 0 56000 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_495
timestamp 1669390400
transform 1 0 56784 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_531
timestamp 1669390400
transform 1 0 60816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_564
timestamp 1669390400
transform 1 0 64512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_570
timestamp 1669390400
transform 1 0 65184 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_578
timestamp 1669390400
transform 1 0 66080 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_582
timestamp 1669390400
transform 1 0 66528 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_613
timestamp 1669390400
transform 1 0 70000 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_623
timestamp 1669390400
transform 1 0 71120 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_627
timestamp 1669390400
transform 1 0 71568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_635
timestamp 1669390400
transform 1 0 72464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_641
timestamp 1669390400
transform 1 0 73136 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_649
timestamp 1669390400
transform 1 0 74032 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_653
timestamp 1669390400
transform 1 0 74480 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_660
timestamp 1669390400
transform 1 0 75264 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_668
timestamp 1669390400
transform 1 0 76160 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_678
timestamp 1669390400
transform 1 0 77280 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_709
timestamp 1669390400
transform 1 0 80752 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_712
timestamp 1669390400
transform 1 0 81088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_742
timestamp 1669390400
transform 1 0 84448 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_773
timestamp 1669390400
transform 1 0 87920 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_777
timestamp 1669390400
transform 1 0 88368 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_783
timestamp 1669390400
transform 1 0 89040 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_787
timestamp 1669390400
transform 1 0 89488 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_789
timestamp 1669390400
transform 1 0 89712 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_840
timestamp 1669390400
transform 1 0 95424 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_848
timestamp 1669390400
transform 1 0 96320 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_854
timestamp 1669390400
transform 1 0 96992 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_862
timestamp 1669390400
transform 1 0 97888 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1669390400
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_424
timestamp 1669390400
transform 1 0 48832 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_440
timestamp 1669390400
transform 1 0 50624 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_447
timestamp 1669390400
transform 1 0 51408 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_455
timestamp 1669390400
transform 1 0 52304 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_459
timestamp 1669390400
transform 1 0 52752 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_479
timestamp 1669390400
transform 1 0 54992 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_510
timestamp 1669390400
transform 1 0 58464 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_514
timestamp 1669390400
transform 1 0 58912 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_530
timestamp 1669390400
transform 1 0 60704 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_534
timestamp 1669390400
transform 1 0 61152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_564
timestamp 1669390400
transform 1 0 64512 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_571
timestamp 1669390400
transform 1 0 65296 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_587
timestamp 1669390400
transform 1 0 67088 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_595
timestamp 1669390400
transform 1 0 67984 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_601
timestamp 1669390400
transform 1 0 68656 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_605
timestamp 1669390400
transform 1 0 69104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_615
timestamp 1669390400
transform 1 0 70224 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_647
timestamp 1669390400
transform 1 0 73808 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_655
timestamp 1669390400
transform 1 0 74704 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_659
timestamp 1669390400
transform 1 0 75152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_662
timestamp 1669390400
transform 1 0 75488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_666
timestamp 1669390400
transform 1 0 75936 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_669
timestamp 1669390400
transform 1 0 76272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1669390400
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_676
timestamp 1669390400
transform 1 0 77056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_679
timestamp 1669390400
transform 1 0 77392 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_687
timestamp 1669390400
transform 1 0 78288 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_689
timestamp 1669390400
transform 1 0 78512 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_696
timestamp 1669390400
transform 1 0 79296 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_704
timestamp 1669390400
transform 1 0 80192 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_710
timestamp 1669390400
transform 1 0 80864 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_718
timestamp 1669390400
transform 1 0 81760 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_735
timestamp 1669390400
transform 1 0 83664 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_739
timestamp 1669390400
transform 1 0 84112 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_741
timestamp 1669390400
transform 1 0 84336 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_744
timestamp 1669390400
transform 1 0 84672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_747
timestamp 1669390400
transform 1 0 85008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_763
timestamp 1669390400
transform 1 0 86800 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_779
timestamp 1669390400
transform 1 0 88592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_785
timestamp 1669390400
transform 1 0 89264 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_787
timestamp 1669390400
transform 1 0 89488 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_793
timestamp 1669390400
transform 1 0 90160 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_795
timestamp 1669390400
transform 1 0 90384 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_801
timestamp 1669390400
transform 1 0 91056 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_805
timestamp 1669390400
transform 1 0 91504 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_811
timestamp 1669390400
transform 1 0 92176 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_815
timestamp 1669390400
transform 1 0 92624 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_818
timestamp 1669390400
transform 1 0 92960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_821
timestamp 1669390400
transform 1 0 93296 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_825
timestamp 1669390400
transform 1 0 93744 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_829
timestamp 1669390400
transform 1 0 94192 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_831
timestamp 1669390400
transform 1 0 94416 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_834
timestamp 1669390400
transform 1 0 94752 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_838
timestamp 1669390400
transform 1 0 95200 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_842
timestamp 1669390400
transform 1 0 95648 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_846
timestamp 1669390400
transform 1 0 96096 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_862
timestamp 1669390400
transform 1 0 97888 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1669390400
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_444
timestamp 1669390400
transform 1 0 51072 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_452
timestamp 1669390400
transform 1 0 51968 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_458
timestamp 1669390400
transform 1 0 52640 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_462
timestamp 1669390400
transform 1 0 53088 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_469
timestamp 1669390400
transform 1 0 53872 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_473
timestamp 1669390400
transform 1 0 54320 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_475
timestamp 1669390400
transform 1 0 54544 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_478
timestamp 1669390400
transform 1 0 54880 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_482
timestamp 1669390400
transform 1 0 55328 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_486
timestamp 1669390400
transform 1 0 55776 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_490
timestamp 1669390400
transform 1 0 56224 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_494
timestamp 1669390400
transform 1 0 56672 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_502
timestamp 1669390400
transform 1 0 57568 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_518
timestamp 1669390400
transform 1 0 59360 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_526
timestamp 1669390400
transform 1 0 60256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_530
timestamp 1669390400
transform 1 0 60704 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_533
timestamp 1669390400
transform 1 0 61040 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_564
timestamp 1669390400
transform 1 0 64512 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_570
timestamp 1669390400
transform 1 0 65184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_576
timestamp 1669390400
transform 1 0 65856 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_580
timestamp 1669390400
transform 1 0 66304 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_582
timestamp 1669390400
transform 1 0 66528 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_612
timestamp 1669390400
transform 1 0 69888 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_616
timestamp 1669390400
transform 1 0 70336 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_620
timestamp 1669390400
transform 1 0 70784 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_628
timestamp 1669390400
transform 1 0 71680 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_631
timestamp 1669390400
transform 1 0 72016 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_635
timestamp 1669390400
transform 1 0 72464 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1669390400
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_641
timestamp 1669390400
transform 1 0 73136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_644
timestamp 1669390400
transform 1 0 73472 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_651
timestamp 1669390400
transform 1 0 74256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_655
timestamp 1669390400
transform 1 0 74704 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_659
timestamp 1669390400
transform 1 0 75152 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_666
timestamp 1669390400
transform 1 0 75936 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_673
timestamp 1669390400
transform 1 0 76720 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_677
timestamp 1669390400
transform 1 0 77168 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_681
timestamp 1669390400
transform 1 0 77616 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_685
timestamp 1669390400
transform 1 0 78064 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_701
timestamp 1669390400
transform 1 0 79856 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_709
timestamp 1669390400
transform 1 0 80752 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_712
timestamp 1669390400
transform 1 0 81088 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_718
timestamp 1669390400
transform 1 0 81760 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_726
timestamp 1669390400
transform 1 0 82656 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_742
timestamp 1669390400
transform 1 0 84448 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_746
timestamp 1669390400
transform 1 0 84896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_749
timestamp 1669390400
transform 1 0 85232 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_780
timestamp 1669390400
transform 1 0 88704 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_783
timestamp 1669390400
transform 1 0 89040 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_816
timestamp 1669390400
transform 1 0 92736 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_823
timestamp 1669390400
transform 1 0 93520 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_827
timestamp 1669390400
transform 1 0 93968 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_831
timestamp 1669390400
transform 1 0 94416 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_835
timestamp 1669390400
transform 1 0 94864 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_839
timestamp 1669390400
transform 1 0 95312 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_843
timestamp 1669390400
transform 1 0 95760 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_847
timestamp 1669390400
transform 1 0 96208 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_851
timestamp 1669390400
transform 1 0 96656 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_854
timestamp 1669390400
transform 1 0 96992 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_862
timestamp 1669390400
transform 1 0 97888 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_385
timestamp 1669390400
transform 1 0 44464 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_424
timestamp 1669390400
transform 1 0 48832 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_426
timestamp 1669390400
transform 1 0 49056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_456
timestamp 1669390400
transform 1 0 52416 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_514
timestamp 1669390400
transform 1 0 58912 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_518
timestamp 1669390400
transform 1 0 59360 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_521
timestamp 1669390400
transform 1 0 59696 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_525
timestamp 1669390400
transform 1 0 60144 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1669390400
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_534
timestamp 1669390400
transform 1 0 61152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_540
timestamp 1669390400
transform 1 0 61824 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_544
timestamp 1669390400
transform 1 0 62272 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_577
timestamp 1669390400
transform 1 0 65968 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_584
timestamp 1669390400
transform 1 0 66752 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_588
timestamp 1669390400
transform 1 0 67200 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_592
timestamp 1669390400
transform 1 0 67648 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_595
timestamp 1669390400
transform 1 0 67984 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1669390400
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_605
timestamp 1669390400
transform 1 0 69104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_611
timestamp 1669390400
transform 1 0 69776 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_618
timestamp 1669390400
transform 1 0 70560 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_622
timestamp 1669390400
transform 1 0 71008 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_626
timestamp 1669390400
transform 1 0 71456 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_630
timestamp 1669390400
transform 1 0 71904 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_636
timestamp 1669390400
transform 1 0 72576 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_667
timestamp 1669390400
transform 1 0 76048 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_671
timestamp 1669390400
transform 1 0 76496 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_673
timestamp 1669390400
transform 1 0 76720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_676
timestamp 1669390400
transform 1 0 77056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_679
timestamp 1669390400
transform 1 0 77392 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_683
timestamp 1669390400
transform 1 0 77840 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_687
timestamp 1669390400
transform 1 0 78288 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_691
timestamp 1669390400
transform 1 0 78736 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_707
timestamp 1669390400
transform 1 0 80528 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_713
timestamp 1669390400
transform 1 0 81200 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_723
timestamp 1669390400
transform 1 0 82320 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_731
timestamp 1669390400
transform 1 0 83216 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_734
timestamp 1669390400
transform 1 0 83552 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_740
timestamp 1669390400
transform 1 0 84224 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_744
timestamp 1669390400
transform 1 0 84672 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_747
timestamp 1669390400
transform 1 0 85008 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_781
timestamp 1669390400
transform 1 0 88816 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_812
timestamp 1669390400
transform 1 0 92288 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_818
timestamp 1669390400
transform 1 0 92960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_825
timestamp 1669390400
transform 1 0 93744 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_832
timestamp 1669390400
transform 1 0 94528 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_836
timestamp 1669390400
transform 1 0 94976 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_840
timestamp 1669390400
transform 1 0 95424 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_844
timestamp 1669390400
transform 1 0 95872 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_850
timestamp 1669390400
transform 1 0 96544 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_854
timestamp 1669390400
transform 1 0 96992 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_858
timestamp 1669390400
transform 1 0 97440 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_421
timestamp 1669390400
transform 1 0 48496 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_430
timestamp 1669390400
transform 1 0 49504 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_460
timestamp 1669390400
transform 1 0 52864 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_467
timestamp 1669390400
transform 1 0 53648 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_474
timestamp 1669390400
transform 1 0 54432 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_481
timestamp 1669390400
transform 1 0 55216 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_485
timestamp 1669390400
transform 1 0 55664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_489
timestamp 1669390400
transform 1 0 56112 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_495
timestamp 1669390400
transform 1 0 56784 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_505
timestamp 1669390400
transform 1 0 57904 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_512
timestamp 1669390400
transform 1 0 58688 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_519
timestamp 1669390400
transform 1 0 59472 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_523
timestamp 1669390400
transform 1 0 59920 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_527
timestamp 1669390400
transform 1 0 60368 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_533
timestamp 1669390400
transform 1 0 61040 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_537
timestamp 1669390400
transform 1 0 61488 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_543
timestamp 1669390400
transform 1 0 62160 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_550
timestamp 1669390400
transform 1 0 62944 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_557
timestamp 1669390400
transform 1 0 63728 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_564
timestamp 1669390400
transform 1 0 64512 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_570
timestamp 1669390400
transform 1 0 65184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_576
timestamp 1669390400
transform 1 0 65856 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_583
timestamp 1669390400
transform 1 0 66640 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_587
timestamp 1669390400
transform 1 0 67088 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_591
timestamp 1669390400
transform 1 0 67536 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_598
timestamp 1669390400
transform 1 0 68320 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_629
timestamp 1669390400
transform 1 0 71792 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_636
timestamp 1669390400
transform 1 0 72576 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1669390400
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_641
timestamp 1669390400
transform 1 0 73136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_644
timestamp 1669390400
transform 1 0 73472 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_675
timestamp 1669390400
transform 1 0 76944 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_709
timestamp 1669390400
transform 1 0 80752 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_712
timestamp 1669390400
transform 1 0 81088 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_714
timestamp 1669390400
transform 1 0 81312 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_744
timestamp 1669390400
transform 1 0 84672 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_775
timestamp 1669390400
transform 1 0 88144 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_777
timestamp 1669390400
transform 1 0 88368 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_780
timestamp 1669390400
transform 1 0 88704 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_783
timestamp 1669390400
transform 1 0 89040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_813
timestamp 1669390400
transform 1 0 92400 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_820
timestamp 1669390400
transform 1 0 93184 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_851
timestamp 1669390400
transform 1 0 96656 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_854
timestamp 1669390400
transform 1 0 96992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_860
timestamp 1669390400
transform 1 0 97664 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_864
timestamp 1669390400
transform 1 0 98112 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_385
timestamp 1669390400
transform 1 0 44464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_424
timestamp 1669390400
transform 1 0 48832 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_428
timestamp 1669390400
transform 1 0 49280 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_430
timestamp 1669390400
transform 1 0 49504 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_469
timestamp 1669390400
transform 1 0 53872 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_476
timestamp 1669390400
transform 1 0 54656 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_483
timestamp 1669390400
transform 1 0 55440 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_514
timestamp 1669390400
transform 1 0 58912 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_522
timestamp 1669390400
transform 1 0 59808 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_526
timestamp 1669390400
transform 1 0 60256 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_528
timestamp 1669390400
transform 1 0 60480 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1669390400
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_534
timestamp 1669390400
transform 1 0 61152 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_538
timestamp 1669390400
transform 1 0 61600 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_590
timestamp 1669390400
transform 1 0 67424 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_594
timestamp 1669390400
transform 1 0 67872 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_596
timestamp 1669390400
transform 1 0 68096 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1669390400
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_605
timestamp 1669390400
transform 1 0 69104 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_607
timestamp 1669390400
transform 1 0 69328 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_658
timestamp 1669390400
transform 1 0 75040 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_666
timestamp 1669390400
transform 1 0 75936 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_670
timestamp 1669390400
transform 1 0 76384 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_676
timestamp 1669390400
transform 1 0 77056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_683
timestamp 1669390400
transform 1 0 77840 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_690
timestamp 1669390400
transform 1 0 78624 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_721
timestamp 1669390400
transform 1 0 82096 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_725
timestamp 1669390400
transform 1 0 82544 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_732
timestamp 1669390400
transform 1 0 83328 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_739
timestamp 1669390400
transform 1 0 84112 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_743
timestamp 1669390400
transform 1 0 84560 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_747
timestamp 1669390400
transform 1 0 85008 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_756
timestamp 1669390400
transform 1 0 86016 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_760
timestamp 1669390400
transform 1 0 86464 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_814
timestamp 1669390400
transform 1 0 92512 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_818
timestamp 1669390400
transform 1 0 92960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_821
timestamp 1669390400
transform 1 0 93296 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_823
timestamp 1669390400
transform 1 0 93520 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_830
timestamp 1669390400
transform 1 0 94304 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_863
timestamp 1669390400
transform 1 0 98000 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_865
timestamp 1669390400
transform 1 0 98224 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_421
timestamp 1669390400
transform 1 0 48496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_444
timestamp 1669390400
transform 1 0 51072 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_448
timestamp 1669390400
transform 1 0 51520 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_478
timestamp 1669390400
transform 1 0 54880 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_486
timestamp 1669390400
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_505
timestamp 1669390400
transform 1 0 57904 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_509
timestamp 1669390400
transform 1 0 58352 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_513
timestamp 1669390400
transform 1 0 58800 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_529
timestamp 1669390400
transform 1 0 60592 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_533
timestamp 1669390400
transform 1 0 61040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_536
timestamp 1669390400
transform 1 0 61376 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1669390400
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_570
timestamp 1669390400
transform 1 0 65184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_576
timestamp 1669390400
transform 1 0 65856 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_583
timestamp 1669390400
transform 1 0 66640 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_587
timestamp 1669390400
transform 1 0 67088 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_591
timestamp 1669390400
transform 1 0 67536 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_593
timestamp 1669390400
transform 1 0 67760 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_600
timestamp 1669390400
transform 1 0 68544 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_604
timestamp 1669390400
transform 1 0 68992 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_612
timestamp 1669390400
transform 1 0 69888 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_620
timestamp 1669390400
transform 1 0 70784 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_628
timestamp 1669390400
transform 1 0 71680 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_635
timestamp 1669390400
transform 1 0 72464 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_641
timestamp 1669390400
transform 1 0 73136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_648
timestamp 1669390400
transform 1 0 73920 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_656
timestamp 1669390400
transform 1 0 74816 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_664
timestamp 1669390400
transform 1 0 75712 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_672
timestamp 1669390400
transform 1 0 76608 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_676
timestamp 1669390400
transform 1 0 77056 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_678
timestamp 1669390400
transform 1 0 77280 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_708
timestamp 1669390400
transform 1 0 80640 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_712
timestamp 1669390400
transform 1 0 81088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_745
timestamp 1669390400
transform 1 0 84784 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_749
timestamp 1669390400
transform 1 0 85232 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_753
timestamp 1669390400
transform 1 0 85680 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_757
timestamp 1669390400
transform 1 0 86128 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_763
timestamp 1669390400
transform 1 0 86800 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_767
timestamp 1669390400
transform 1 0 87248 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_773
timestamp 1669390400
transform 1 0 87920 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_780
timestamp 1669390400
transform 1 0 88704 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_783
timestamp 1669390400
transform 1 0 89040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_789
timestamp 1669390400
transform 1 0 89712 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_796
timestamp 1669390400
transform 1 0 90496 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_800
timestamp 1669390400
transform 1 0 90944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_830
timestamp 1669390400
transform 1 0 94304 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_837
timestamp 1669390400
transform 1 0 95088 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_844
timestamp 1669390400
transform 1 0 95872 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_851
timestamp 1669390400
transform 1 0 96656 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_854
timestamp 1669390400
transform 1 0 96992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_860
timestamp 1669390400
transform 1 0 97664 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_864
timestamp 1669390400
transform 1 0 98112 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_424
timestamp 1669390400
transform 1 0 48832 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_440
timestamp 1669390400
transform 1 0 50624 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_442
timestamp 1669390400
transform 1 0 50848 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_445
timestamp 1669390400
transform 1 0 51184 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_453
timestamp 1669390400
transform 1 0 52080 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_469
timestamp 1669390400
transform 1 0 53872 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_476
timestamp 1669390400
transform 1 0 54656 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_478
timestamp 1669390400
transform 1 0 54880 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_511
timestamp 1669390400
transform 1 0 58576 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_515
timestamp 1669390400
transform 1 0 59024 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_519
timestamp 1669390400
transform 1 0 59472 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_523
timestamp 1669390400
transform 1 0 59920 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_527
timestamp 1669390400
transform 1 0 60368 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_531
timestamp 1669390400
transform 1 0 60816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_534
timestamp 1669390400
transform 1 0 61152 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_538
timestamp 1669390400
transform 1 0 61600 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_568
timestamp 1669390400
transform 1 0 64960 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_575
timestamp 1669390400
transform 1 0 65744 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_579
timestamp 1669390400
transform 1 0 66192 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_583
timestamp 1669390400
transform 1 0 66640 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_599
timestamp 1669390400
transform 1 0 68432 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_605
timestamp 1669390400
transform 1 0 69104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_608
timestamp 1669390400
transform 1 0 69440 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_615
timestamp 1669390400
transform 1 0 70224 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_619
timestamp 1669390400
transform 1 0 70672 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_650
timestamp 1669390400
transform 1 0 74144 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_654
timestamp 1669390400
transform 1 0 74592 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_661
timestamp 1669390400
transform 1 0 75376 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_663
timestamp 1669390400
transform 1 0 75600 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_670
timestamp 1669390400
transform 1 0 76384 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_676
timestamp 1669390400
transform 1 0 77056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_679
timestamp 1669390400
transform 1 0 77392 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_683
timestamp 1669390400
transform 1 0 77840 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_734
timestamp 1669390400
transform 1 0 83552 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_738
timestamp 1669390400
transform 1 0 84000 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_742
timestamp 1669390400
transform 1 0 84448 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_744
timestamp 1669390400
transform 1 0 84672 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_747
timestamp 1669390400
transform 1 0 85008 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_751
timestamp 1669390400
transform 1 0 85456 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_755
timestamp 1669390400
transform 1 0 85904 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_763
timestamp 1669390400
transform 1 0 86800 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_765
timestamp 1669390400
transform 1 0 87024 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_768
timestamp 1669390400
transform 1 0 87360 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_776
timestamp 1669390400
transform 1 0 88256 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_780
timestamp 1669390400
transform 1 0 88704 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_783
timestamp 1669390400
transform 1 0 89040 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_787
timestamp 1669390400
transform 1 0 89488 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_794
timestamp 1669390400
transform 1 0 90272 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_803
timestamp 1669390400
transform 1 0 91280 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_810
timestamp 1669390400
transform 1 0 92064 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_814
timestamp 1669390400
transform 1 0 92512 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_818
timestamp 1669390400
transform 1 0 92960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_824
timestamp 1669390400
transform 1 0 93632 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_831
timestamp 1669390400
transform 1 0 94416 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_833
timestamp 1669390400
transform 1 0 94640 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_863
timestamp 1669390400
transform 1 0 98000 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_865
timestamp 1669390400
transform 1 0 98224 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_421
timestamp 1669390400
transform 1 0 48496 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_460
timestamp 1669390400
transform 1 0 52864 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_464
timestamp 1669390400
transform 1 0 53312 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_474
timestamp 1669390400
transform 1 0 54432 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_478
timestamp 1669390400
transform 1 0 54880 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_482
timestamp 1669390400
transform 1 0 55328 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_486
timestamp 1669390400
transform 1 0 55776 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_490
timestamp 1669390400
transform 1 0 56224 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_494
timestamp 1669390400
transform 1 0 56672 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_502
timestamp 1669390400
transform 1 0 57568 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_536
timestamp 1669390400
transform 1 0 61376 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_540
timestamp 1669390400
transform 1 0 61824 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_544
timestamp 1669390400
transform 1 0 62272 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_548
timestamp 1669390400
transform 1 0 62720 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_552
timestamp 1669390400
transform 1 0 63168 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_556
timestamp 1669390400
transform 1 0 63616 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_562
timestamp 1669390400
transform 1 0 64288 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_566
timestamp 1669390400
transform 1 0 64736 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_570
timestamp 1669390400
transform 1 0 65184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_573
timestamp 1669390400
transform 1 0 65520 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_581
timestamp 1669390400
transform 1 0 66416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_585
timestamp 1669390400
transform 1 0 66864 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_616
timestamp 1669390400
transform 1 0 70336 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_620
timestamp 1669390400
transform 1 0 70784 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_624
timestamp 1669390400
transform 1 0 71232 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_630
timestamp 1669390400
transform 1 0 71904 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1669390400
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_641
timestamp 1669390400
transform 1 0 73136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_647
timestamp 1669390400
transform 1 0 73808 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_651
timestamp 1669390400
transform 1 0 74256 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_655
timestamp 1669390400
transform 1 0 74704 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_659
timestamp 1669390400
transform 1 0 75152 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_667
timestamp 1669390400
transform 1 0 76048 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_671
timestamp 1669390400
transform 1 0 76496 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_677
timestamp 1669390400
transform 1 0 77168 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_681
timestamp 1669390400
transform 1 0 77616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_690
timestamp 1669390400
transform 1 0 78624 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_692
timestamp 1669390400
transform 1 0 78848 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_698
timestamp 1669390400
transform 1 0 79520 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_705
timestamp 1669390400
transform 1 0 80304 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_709
timestamp 1669390400
transform 1 0 80752 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_712
timestamp 1669390400
transform 1 0 81088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_718
timestamp 1669390400
transform 1 0 81760 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_722
timestamp 1669390400
transform 1 0 82208 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_726
timestamp 1669390400
transform 1 0 82656 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_742
timestamp 1669390400
transform 1 0 84448 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_750
timestamp 1669390400
transform 1 0 85344 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_752
timestamp 1669390400
transform 1 0 85568 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_755
timestamp 1669390400
transform 1 0 85904 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_771
timestamp 1669390400
transform 1 0 87696 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_779
timestamp 1669390400
transform 1 0 88592 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_783
timestamp 1669390400
transform 1 0 89040 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_789
timestamp 1669390400
transform 1 0 89712 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_793
timestamp 1669390400
transform 1 0 90160 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_797
timestamp 1669390400
transform 1 0 90608 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_851
timestamp 1669390400
transform 1 0 96656 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_854
timestamp 1669390400
transform 1 0 96992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_860
timestamp 1669390400
transform 1 0 97664 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_864
timestamp 1669390400
transform 1 0 98112 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_424
timestamp 1669390400
transform 1 0 48832 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_426
timestamp 1669390400
transform 1 0 49056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_433
timestamp 1669390400
transform 1 0 49840 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_449
timestamp 1669390400
transform 1 0 51632 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_457
timestamp 1669390400
transform 1 0 52528 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_466
timestamp 1669390400
transform 1 0 53536 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_470
timestamp 1669390400
transform 1 0 53984 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_506
timestamp 1669390400
transform 1 0 58016 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_510
timestamp 1669390400
transform 1 0 58464 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_514
timestamp 1669390400
transform 1 0 58912 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_530
timestamp 1669390400
transform 1 0 60704 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_534
timestamp 1669390400
transform 1 0 61152 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_542
timestamp 1669390400
transform 1 0 62048 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_545
timestamp 1669390400
transform 1 0 62384 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_549
timestamp 1669390400
transform 1 0 62832 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_565
timestamp 1669390400
transform 1 0 64624 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_573
timestamp 1669390400
transform 1 0 65520 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_577
timestamp 1669390400
transform 1 0 65968 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_581
timestamp 1669390400
transform 1 0 66416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_590
timestamp 1669390400
transform 1 0 67424 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_597
timestamp 1669390400
transform 1 0 68208 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_601
timestamp 1669390400
transform 1 0 68656 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_605
timestamp 1669390400
transform 1 0 69104 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_609
timestamp 1669390400
transform 1 0 69552 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_642
timestamp 1669390400
transform 1 0 73248 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_646
timestamp 1669390400
transform 1 0 73696 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_650
timestamp 1669390400
transform 1 0 74144 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_660
timestamp 1669390400
transform 1 0 75264 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_662
timestamp 1669390400
transform 1 0 75488 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_671
timestamp 1669390400
transform 1 0 76496 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_673
timestamp 1669390400
transform 1 0 76720 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_676
timestamp 1669390400
transform 1 0 77056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_679
timestamp 1669390400
transform 1 0 77392 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_683
timestamp 1669390400
transform 1 0 77840 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_693
timestamp 1669390400
transform 1 0 78960 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_725
timestamp 1669390400
transform 1 0 82544 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_741
timestamp 1669390400
transform 1 0 84336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_747
timestamp 1669390400
transform 1 0 85008 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_753
timestamp 1669390400
transform 1 0 85680 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_787
timestamp 1669390400
transform 1 0 89488 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_795
timestamp 1669390400
transform 1 0 90384 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_799
timestamp 1669390400
transform 1 0 90832 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_806
timestamp 1669390400
transform 1 0 91616 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_810
timestamp 1669390400
transform 1 0 92064 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_814
timestamp 1669390400
transform 1 0 92512 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_818
timestamp 1669390400
transform 1 0 92960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_824
timestamp 1669390400
transform 1 0 93632 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_831
timestamp 1669390400
transform 1 0 94416 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_862
timestamp 1669390400
transform 1 0 97888 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_421
timestamp 1669390400
transform 1 0 48496 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_458
timestamp 1669390400
transform 1 0 52640 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_462
timestamp 1669390400
transform 1 0 53088 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_494
timestamp 1669390400
transform 1 0 56672 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_531
timestamp 1669390400
transform 1 0 60816 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_533
timestamp 1669390400
transform 1 0 61040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_536
timestamp 1669390400
transform 1 0 61376 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_543
timestamp 1669390400
transform 1 0 62160 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_550
timestamp 1669390400
transform 1 0 62944 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_557
timestamp 1669390400
transform 1 0 63728 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_561
timestamp 1669390400
transform 1 0 64176 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_565
timestamp 1669390400
transform 1 0 64624 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_567
timestamp 1669390400
transform 1 0 64848 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_570
timestamp 1669390400
transform 1 0 65184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_573
timestamp 1669390400
transform 1 0 65520 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_577
timestamp 1669390400
transform 1 0 65968 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_610
timestamp 1669390400
transform 1 0 69664 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_614
timestamp 1669390400
transform 1 0 70112 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_617
timestamp 1669390400
transform 1 0 70448 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_625
timestamp 1669390400
transform 1 0 71344 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_635
timestamp 1669390400
transform 1 0 72464 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_641
timestamp 1669390400
transform 1 0 73136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_650
timestamp 1669390400
transform 1 0 74144 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_654
timestamp 1669390400
transform 1 0 74592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_658
timestamp 1669390400
transform 1 0 75040 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_662
timestamp 1669390400
transform 1 0 75488 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_666
timestamp 1669390400
transform 1 0 75936 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_674
timestamp 1669390400
transform 1 0 76832 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_678
timestamp 1669390400
transform 1 0 77280 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_680
timestamp 1669390400
transform 1 0 77504 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_683
timestamp 1669390400
transform 1 0 77840 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_685
timestamp 1669390400
transform 1 0 78064 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_691
timestamp 1669390400
transform 1 0 78736 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_695
timestamp 1669390400
transform 1 0 79184 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_699
timestamp 1669390400
transform 1 0 79632 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_707
timestamp 1669390400
transform 1 0 80528 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_709
timestamp 1669390400
transform 1 0 80752 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_712
timestamp 1669390400
transform 1 0 81088 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_730
timestamp 1669390400
transform 1 0 83104 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_746
timestamp 1669390400
transform 1 0 84896 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_777
timestamp 1669390400
transform 1 0 88368 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_783
timestamp 1669390400
transform 1 0 89040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_789
timestamp 1669390400
transform 1 0 89712 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_793
timestamp 1669390400
transform 1 0 90160 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_797
timestamp 1669390400
transform 1 0 90608 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_801
timestamp 1669390400
transform 1 0 91056 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_809
timestamp 1669390400
transform 1 0 91952 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_812
timestamp 1669390400
transform 1 0 92288 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_814
timestamp 1669390400
transform 1 0 92512 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_817
timestamp 1669390400
transform 1 0 92848 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_821
timestamp 1669390400
transform 1 0 93296 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_825
timestamp 1669390400
transform 1 0 93744 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_829
timestamp 1669390400
transform 1 0 94192 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_836
timestamp 1669390400
transform 1 0 94976 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_843
timestamp 1669390400
transform 1 0 95760 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_850
timestamp 1669390400
transform 1 0 96544 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_854
timestamp 1669390400
transform 1 0 96992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_857
timestamp 1669390400
transform 1 0 97328 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_861
timestamp 1669390400
transform 1 0 97776 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_865
timestamp 1669390400
transform 1 0 98224 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_408
timestamp 1669390400
transform 1 0 47040 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_412
timestamp 1669390400
transform 1 0 47488 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_420
timestamp 1669390400
transform 1 0 48384 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_451
timestamp 1669390400
transform 1 0 51856 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_455
timestamp 1669390400
transform 1 0 52304 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_459
timestamp 1669390400
transform 1 0 52752 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_479
timestamp 1669390400
transform 1 0 54992 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_487
timestamp 1669390400
transform 1 0 55888 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_489
timestamp 1669390400
transform 1 0 56112 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_499
timestamp 1669390400
transform 1 0 57232 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_503
timestamp 1669390400
transform 1 0 57680 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_519
timestamp 1669390400
transform 1 0 59472 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_523
timestamp 1669390400
transform 1 0 59920 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_525
timestamp 1669390400
transform 1 0 60144 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_528
timestamp 1669390400
transform 1 0 60480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_534
timestamp 1669390400
transform 1 0 61152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_564
timestamp 1669390400
transform 1 0 64512 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_568
timestamp 1669390400
transform 1 0 64960 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_570
timestamp 1669390400
transform 1 0 65184 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_576
timestamp 1669390400
transform 1 0 65856 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_580
timestamp 1669390400
transform 1 0 66304 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_584
timestamp 1669390400
transform 1 0 66752 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_588
timestamp 1669390400
transform 1 0 67200 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_595
timestamp 1669390400
transform 1 0 67984 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1669390400
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_605
timestamp 1669390400
transform 1 0 69104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_611
timestamp 1669390400
transform 1 0 69776 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_618
timestamp 1669390400
transform 1 0 70560 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_622
timestamp 1669390400
transform 1 0 71008 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_626
timestamp 1669390400
transform 1 0 71456 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_634
timestamp 1669390400
transform 1 0 72352 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_637
timestamp 1669390400
transform 1 0 72688 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_639
timestamp 1669390400
transform 1 0 72912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_642
timestamp 1669390400
transform 1 0 73248 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_646
timestamp 1669390400
transform 1 0 73696 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_656
timestamp 1669390400
transform 1 0 74816 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_666
timestamp 1669390400
transform 1 0 75936 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_673
timestamp 1669390400
transform 1 0 76720 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_676
timestamp 1669390400
transform 1 0 77056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_706
timestamp 1669390400
transform 1 0 80416 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_710
timestamp 1669390400
transform 1 0 80864 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_718
timestamp 1669390400
transform 1 0 81760 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_722
timestamp 1669390400
transform 1 0 82208 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_725
timestamp 1669390400
transform 1 0 82544 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_742
timestamp 1669390400
transform 1 0 84448 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_744
timestamp 1669390400
transform 1 0 84672 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_747
timestamp 1669390400
transform 1 0 85008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_750
timestamp 1669390400
transform 1 0 85344 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_758
timestamp 1669390400
transform 1 0 86240 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_761
timestamp 1669390400
transform 1 0 86576 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_768
timestamp 1669390400
transform 1 0 87360 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_770
timestamp 1669390400
transform 1 0 87584 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_800
timestamp 1669390400
transform 1 0 90944 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_804
timestamp 1669390400
transform 1 0 91392 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_808
timestamp 1669390400
transform 1 0 91840 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_810
timestamp 1669390400
transform 1 0 92064 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_813
timestamp 1669390400
transform 1 0 92400 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_815
timestamp 1669390400
transform 1 0 92624 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_818
timestamp 1669390400
transform 1 0 92960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_821
timestamp 1669390400
transform 1 0 93296 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_825
timestamp 1669390400
transform 1 0 93744 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_829
timestamp 1669390400
transform 1 0 94192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_862
timestamp 1669390400
transform 1 0 97888 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_389
timestamp 1669390400
transform 1 0 44912 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_405
timestamp 1669390400
transform 1 0 46704 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_413
timestamp 1669390400
transform 1 0 47600 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_417
timestamp 1669390400
transform 1 0 48048 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_430
timestamp 1669390400
transform 1 0 49504 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_446
timestamp 1669390400
transform 1 0 51296 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_463
timestamp 1669390400
transform 1 0 53200 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_467
timestamp 1669390400
transform 1 0 53648 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_471
timestamp 1669390400
transform 1 0 54096 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_475
timestamp 1669390400
transform 1 0 54544 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_481
timestamp 1669390400
transform 1 0 55216 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_488
timestamp 1669390400
transform 1 0 56000 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_495
timestamp 1669390400
transform 1 0 56784 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_502
timestamp 1669390400
transform 1 0 57568 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_506
timestamp 1669390400
transform 1 0 58016 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_514
timestamp 1669390400
transform 1 0 58912 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_516
timestamp 1669390400
transform 1 0 59136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_519
timestamp 1669390400
transform 1 0 59472 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_526
timestamp 1669390400
transform 1 0 60256 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_557
timestamp 1669390400
transform 1 0 63728 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_564
timestamp 1669390400
transform 1 0 64512 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_570
timestamp 1669390400
transform 1 0 65184 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_572
timestamp 1669390400
transform 1 0 65408 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_602
timestamp 1669390400
transform 1 0 68768 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_610
timestamp 1669390400
transform 1 0 69664 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_614
timestamp 1669390400
transform 1 0 70112 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_622
timestamp 1669390400
transform 1 0 71008 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_625
timestamp 1669390400
transform 1 0 71344 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_627
timestamp 1669390400
transform 1 0 71568 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_630
timestamp 1669390400
transform 1 0 71904 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_634
timestamp 1669390400
transform 1 0 72352 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1669390400
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_641
timestamp 1669390400
transform 1 0 73136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_654
timestamp 1669390400
transform 1 0 74592 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_664
timestamp 1669390400
transform 1 0 75712 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_668
timestamp 1669390400
transform 1 0 76160 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_675
timestamp 1669390400
transform 1 0 76944 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_679
timestamp 1669390400
transform 1 0 77392 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_709
timestamp 1669390400
transform 1 0 80752 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_712
timestamp 1669390400
transform 1 0 81088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_715
timestamp 1669390400
transform 1 0 81424 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_746
timestamp 1669390400
transform 1 0 84896 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_754
timestamp 1669390400
transform 1 0 85792 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_758
timestamp 1669390400
transform 1 0 86240 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_762
timestamp 1669390400
transform 1 0 86688 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_765
timestamp 1669390400
transform 1 0 87024 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_772
timestamp 1669390400
transform 1 0 87808 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_779
timestamp 1669390400
transform 1 0 88592 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_783
timestamp 1669390400
transform 1 0 89040 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_790
timestamp 1669390400
transform 1 0 89824 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_797
timestamp 1669390400
transform 1 0 90608 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_804
timestamp 1669390400
transform 1 0 91392 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_808
timestamp 1669390400
transform 1 0 91840 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_812
timestamp 1669390400
transform 1 0 92288 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_814
timestamp 1669390400
transform 1 0 92512 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_820
timestamp 1669390400
transform 1 0 93184 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_827
timestamp 1669390400
transform 1 0 93968 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_834
timestamp 1669390400
transform 1 0 94752 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_838
timestamp 1669390400
transform 1 0 95200 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_846
timestamp 1669390400
transform 1 0 96096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_850
timestamp 1669390400
transform 1 0 96544 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_854
timestamp 1669390400
transform 1 0 96992 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_864
timestamp 1669390400
transform 1 0 98112 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1669390400
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_408
timestamp 1669390400
transform 1 0 47040 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_416
timestamp 1669390400
transform 1 0 47936 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_447
timestamp 1669390400
transform 1 0 51408 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_455
timestamp 1669390400
transform 1 0 52304 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_459
timestamp 1669390400
transform 1 0 52752 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_465
timestamp 1669390400
transform 1 0 53424 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_495
timestamp 1669390400
transform 1 0 56784 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_499
timestamp 1669390400
transform 1 0 57232 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_515
timestamp 1669390400
transform 1 0 59024 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_523
timestamp 1669390400
transform 1 0 59920 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_527
timestamp 1669390400
transform 1 0 60368 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1669390400
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_534
timestamp 1669390400
transform 1 0 61152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_537
timestamp 1669390400
transform 1 0 61488 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_541
timestamp 1669390400
transform 1 0 61936 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_547
timestamp 1669390400
transform 1 0 62608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_551
timestamp 1669390400
transform 1 0 63056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1669390400
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_605
timestamp 1669390400
transform 1 0 69104 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_613
timestamp 1669390400
transform 1 0 70000 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_623
timestamp 1669390400
transform 1 0 71120 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_627
timestamp 1669390400
transform 1 0 71568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_634
timestamp 1669390400
transform 1 0 72352 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_673
timestamp 1669390400
transform 1 0 76720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_676
timestamp 1669390400
transform 1 0 77056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_679
timestamp 1669390400
transform 1 0 77392 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_689
timestamp 1669390400
transform 1 0 78512 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_696
timestamp 1669390400
transform 1 0 79296 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_698
timestamp 1669390400
transform 1 0 79520 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_728
timestamp 1669390400
transform 1 0 82880 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_736
timestamp 1669390400
transform 1 0 83776 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_744
timestamp 1669390400
transform 1 0 84672 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_747
timestamp 1669390400
transform 1 0 85008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_777
timestamp 1669390400
transform 1 0 88368 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_810
timestamp 1669390400
transform 1 0 92064 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_814
timestamp 1669390400
transform 1 0 92512 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_818
timestamp 1669390400
transform 1 0 92960 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_851
timestamp 1669390400
transform 1 0 96656 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_855
timestamp 1669390400
transform 1 0 97104 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_863
timestamp 1669390400
transform 1 0 98000 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_865
timestamp 1669390400
transform 1 0 98224 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_66
timestamp 1669390400
transform 1 0 8736 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1669390400
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1669390400
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1669390400
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_208
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1669390400
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1669390400
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_350
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_421
timestamp 1669390400
transform 1 0 48496 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1669390400
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_428
timestamp 1669390400
transform 1 0 49280 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_436
timestamp 1669390400
transform 1 0 50176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_442
timestamp 1669390400
transform 1 0 50848 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_494
timestamp 1669390400
transform 1 0 56672 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1669390400
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_499
timestamp 1669390400
transform 1 0 57232 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_505
timestamp 1669390400
transform 1 0 57904 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_509
timestamp 1669390400
transform 1 0 58352 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_525
timestamp 1669390400
transform 1 0 60144 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_529
timestamp 1669390400
transform 1 0 60592 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_535
timestamp 1669390400
transform 1 0 61264 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_566
timestamp 1669390400
transform 1 0 64736 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_570
timestamp 1669390400
transform 1 0 65184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_576
timestamp 1669390400
transform 1 0 65856 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_580
timestamp 1669390400
transform 1 0 66304 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_593
timestamp 1669390400
transform 1 0 67760 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_600
timestamp 1669390400
transform 1 0 68544 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_604
timestamp 1669390400
transform 1 0 68992 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_620
timestamp 1669390400
transform 1 0 70784 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_623
timestamp 1669390400
transform 1 0 71120 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_627
timestamp 1669390400
transform 1 0 71568 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_631
timestamp 1669390400
transform 1 0 72016 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1669390400
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_641
timestamp 1669390400
transform 1 0 73136 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_650
timestamp 1669390400
transform 1 0 74144 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_658
timestamp 1669390400
transform 1 0 75040 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_666
timestamp 1669390400
transform 1 0 75936 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_674
timestamp 1669390400
transform 1 0 76832 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_681
timestamp 1669390400
transform 1 0 77616 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_685
timestamp 1669390400
transform 1 0 78064 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_689
timestamp 1669390400
transform 1 0 78512 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_695
timestamp 1669390400
transform 1 0 79184 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_699
timestamp 1669390400
transform 1 0 79632 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_707
timestamp 1669390400
transform 1 0 80528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_709
timestamp 1669390400
transform 1 0 80752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_712
timestamp 1669390400
transform 1 0 81088 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_766
timestamp 1669390400
transform 1 0 87136 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_770
timestamp 1669390400
transform 1 0 87584 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_774
timestamp 1669390400
transform 1 0 88032 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_780
timestamp 1669390400
transform 1 0 88704 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_783
timestamp 1669390400
transform 1 0 89040 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_792
timestamp 1669390400
transform 1 0 90048 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_799
timestamp 1669390400
transform 1 0 90832 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_851
timestamp 1669390400
transform 1 0 96656 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_854
timestamp 1669390400
transform 1 0 96992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_857
timestamp 1669390400
transform 1 0 97328 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_865
timestamp 1669390400
transform 1 0 98224 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1669390400
transform 1 0 5152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1669390400
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_101
timestamp 1669390400
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1669390400
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1669390400
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_172
timestamp 1669390400
transform 1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1669390400
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1669390400
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_243
timestamp 1669390400
transform 1 0 28560 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1669390400
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1669390400
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_314
timestamp 1669390400
transform 1 0 36512 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1669390400
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1669390400
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_385
timestamp 1669390400
transform 1 0 44464 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1669390400
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_392
timestamp 1669390400
transform 1 0 45248 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_408
timestamp 1669390400
transform 1 0 47040 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_416
timestamp 1669390400
transform 1 0 47936 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_447
timestamp 1669390400
transform 1 0 51408 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_451
timestamp 1669390400
transform 1 0 51856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_455
timestamp 1669390400
transform 1 0 52304 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_457
timestamp 1669390400
transform 1 0 52528 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1669390400
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_463
timestamp 1669390400
transform 1 0 53200 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_494
timestamp 1669390400
transform 1 0 56672 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_503
timestamp 1669390400
transform 1 0 57680 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_510
timestamp 1669390400
transform 1 0 58464 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_514
timestamp 1669390400
transform 1 0 58912 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_68_518
timestamp 1669390400
transform 1 0 59360 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_526
timestamp 1669390400
transform 1 0 60256 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_530
timestamp 1669390400
transform 1 0 60704 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_534
timestamp 1669390400
transform 1 0 61152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_564
timestamp 1669390400
transform 1 0 64512 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_568
timestamp 1669390400
transform 1 0 64960 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_572
timestamp 1669390400
transform 1 0 65408 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_588
timestamp 1669390400
transform 1 0 67200 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_592
timestamp 1669390400
transform 1 0 67648 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1669390400
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_605
timestamp 1669390400
transform 1 0 69104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_612
timestamp 1669390400
transform 1 0 69888 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_616
timestamp 1669390400
transform 1 0 70336 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_620
timestamp 1669390400
transform 1 0 70784 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_624
timestamp 1669390400
transform 1 0 71232 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_632
timestamp 1669390400
transform 1 0 72128 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_642
timestamp 1669390400
transform 1 0 73248 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_654
timestamp 1669390400
transform 1 0 74592 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_662
timestamp 1669390400
transform 1 0 75488 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_668
timestamp 1669390400
transform 1 0 76160 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_672
timestamp 1669390400
transform 1 0 76608 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_676
timestamp 1669390400
transform 1 0 77056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_679
timestamp 1669390400
transform 1 0 77392 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_683
timestamp 1669390400
transform 1 0 77840 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_714
timestamp 1669390400
transform 1 0 81312 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_721
timestamp 1669390400
transform 1 0 82096 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_727
timestamp 1669390400
transform 1 0 82768 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_744
timestamp 1669390400
transform 1 0 84672 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_747
timestamp 1669390400
transform 1 0 85008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_750
timestamp 1669390400
transform 1 0 85344 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_766
timestamp 1669390400
transform 1 0 87136 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_770
timestamp 1669390400
transform 1 0 87584 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_772
timestamp 1669390400
transform 1 0 87808 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_775
timestamp 1669390400
transform 1 0 88144 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_782
timestamp 1669390400
transform 1 0 88928 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_813
timestamp 1669390400
transform 1 0 92400 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_815
timestamp 1669390400
transform 1 0 92624 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_818
timestamp 1669390400
transform 1 0 92960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_824
timestamp 1669390400
transform 1 0 93632 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_857
timestamp 1669390400
transform 1 0 97328 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_861
timestamp 1669390400
transform 1 0 97776 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_865
timestamp 1669390400
transform 1 0 98224 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_66
timestamp 1669390400
transform 1 0 8736 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1669390400
transform 1 0 9184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1669390400
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_137
timestamp 1669390400
transform 1 0 16688 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1669390400
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1669390400
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_208
timestamp 1669390400
transform 1 0 24640 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1669390400
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1669390400
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_279
timestamp 1669390400
transform 1 0 32592 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1669390400
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1669390400
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_350
timestamp 1669390400
transform 1 0 40544 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1669390400
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_421
timestamp 1669390400
transform 1 0 48496 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1669390400
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_428
timestamp 1669390400
transform 1 0 49280 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_444
timestamp 1669390400
transform 1 0 51072 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_452
timestamp 1669390400
transform 1 0 51968 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_456
timestamp 1669390400
transform 1 0 52416 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_465
timestamp 1669390400
transform 1 0 53424 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1669390400
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_499
timestamp 1669390400
transform 1 0 57232 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_505
timestamp 1669390400
transform 1 0 57904 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_563
timestamp 1669390400
transform 1 0 64400 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1669390400
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_570
timestamp 1669390400
transform 1 0 65184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_576
timestamp 1669390400
transform 1 0 65856 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_580
timestamp 1669390400
transform 1 0 66304 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_584
timestamp 1669390400
transform 1 0 66752 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_593
timestamp 1669390400
transform 1 0 67760 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_597
timestamp 1669390400
transform 1 0 68208 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_601
timestamp 1669390400
transform 1 0 68656 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_604
timestamp 1669390400
transform 1 0 68992 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_610
timestamp 1669390400
transform 1 0 69664 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_614
timestamp 1669390400
transform 1 0 70112 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_618
timestamp 1669390400
transform 1 0 70560 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_622
timestamp 1669390400
transform 1 0 71008 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_634
timestamp 1669390400
transform 1 0 72352 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1669390400
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_641
timestamp 1669390400
transform 1 0 73136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_647
timestamp 1669390400
transform 1 0 73808 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_660
timestamp 1669390400
transform 1 0 75264 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_671
timestamp 1669390400
transform 1 0 76496 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_677
timestamp 1669390400
transform 1 0 77168 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_681
timestamp 1669390400
transform 1 0 77616 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_685
timestamp 1669390400
transform 1 0 78064 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_687
timestamp 1669390400
transform 1 0 78288 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_694
timestamp 1669390400
transform 1 0 79072 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_701
timestamp 1669390400
transform 1 0 79856 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_703
timestamp 1669390400
transform 1 0 80080 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_709
timestamp 1669390400
transform 1 0 80752 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_712
timestamp 1669390400
transform 1 0 81088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_718
timestamp 1669390400
transform 1 0 81760 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_722
timestamp 1669390400
transform 1 0 82208 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_726
timestamp 1669390400
transform 1 0 82656 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_730
timestamp 1669390400
transform 1 0 83104 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_766
timestamp 1669390400
transform 1 0 87136 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_69_770
timestamp 1669390400
transform 1 0 87584 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_774
timestamp 1669390400
transform 1 0 88032 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_780
timestamp 1669390400
transform 1 0 88704 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_783
timestamp 1669390400
transform 1 0 89040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_813
timestamp 1669390400
transform 1 0 92400 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_820
timestamp 1669390400
transform 1 0 93184 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_851
timestamp 1669390400
transform 1 0 96656 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_854
timestamp 1669390400
transform 1 0 96992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_860
timestamp 1669390400
transform 1 0 97664 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_864
timestamp 1669390400
transform 1 0 98112 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_34
timestamp 1669390400
transform 1 0 5152 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1669390400
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_101
timestamp 1669390400
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1669390400
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1669390400
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_172
timestamp 1669390400
transform 1 0 20608 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1669390400
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1669390400
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_243
timestamp 1669390400
transform 1 0 28560 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1669390400
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1669390400
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_314
timestamp 1669390400
transform 1 0 36512 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1669390400
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1669390400
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_385
timestamp 1669390400
transform 1 0 44464 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1669390400
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_392
timestamp 1669390400
transform 1 0 45248 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_408
timestamp 1669390400
transform 1 0 47040 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_412
timestamp 1669390400
transform 1 0 47488 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_414
timestamp 1669390400
transform 1 0 47712 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_417
timestamp 1669390400
transform 1 0 48048 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_425
timestamp 1669390400
transform 1 0 48944 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_442
timestamp 1669390400
transform 1 0 50848 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_446
timestamp 1669390400
transform 1 0 51296 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_450
timestamp 1669390400
transform 1 0 51744 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_454
timestamp 1669390400
transform 1 0 52192 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1669390400
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_463
timestamp 1669390400
transform 1 0 53200 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_467
timestamp 1669390400
transform 1 0 53648 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_471
timestamp 1669390400
transform 1 0 54096 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_477
timestamp 1669390400
transform 1 0 54768 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_508
timestamp 1669390400
transform 1 0 58240 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_512
timestamp 1669390400
transform 1 0 58688 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_520
timestamp 1669390400
transform 1 0 59584 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_524
timestamp 1669390400
transform 1 0 60032 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1669390400
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_534
timestamp 1669390400
transform 1 0 61152 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_564
timestamp 1669390400
transform 1 0 64512 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_571
timestamp 1669390400
transform 1 0 65296 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_578
timestamp 1669390400
transform 1 0 66080 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_582
timestamp 1669390400
transform 1 0 66528 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_586
timestamp 1669390400
transform 1 0 66976 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_594
timestamp 1669390400
transform 1 0 67872 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_598
timestamp 1669390400
transform 1 0 68320 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1669390400
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_605
timestamp 1669390400
transform 1 0 69104 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_609
timestamp 1669390400
transform 1 0 69552 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_613
timestamp 1669390400
transform 1 0 70000 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_617
timestamp 1669390400
transform 1 0 70448 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_625
timestamp 1669390400
transform 1 0 71344 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_636
timestamp 1669390400
transform 1 0 72576 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_640
timestamp 1669390400
transform 1 0 73024 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_658
timestamp 1669390400
transform 1 0 75040 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_669
timestamp 1669390400
transform 1 0 76272 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_673
timestamp 1669390400
transform 1 0 76720 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_676
timestamp 1669390400
transform 1 0 77056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_683
timestamp 1669390400
transform 1 0 77840 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_690
timestamp 1669390400
transform 1 0 78624 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_694
timestamp 1669390400
transform 1 0 79072 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_698
timestamp 1669390400
transform 1 0 79520 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_702
timestamp 1669390400
transform 1 0 79968 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_706
timestamp 1669390400
transform 1 0 80416 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_710
timestamp 1669390400
transform 1 0 80864 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_714
timestamp 1669390400
transform 1 0 81312 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_718
timestamp 1669390400
transform 1 0 81760 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_722
timestamp 1669390400
transform 1 0 82208 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_732
timestamp 1669390400
transform 1 0 83328 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_736
timestamp 1669390400
transform 1 0 83776 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_740
timestamp 1669390400
transform 1 0 84224 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_744
timestamp 1669390400
transform 1 0 84672 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_747
timestamp 1669390400
transform 1 0 85008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_750
timestamp 1669390400
transform 1 0 85344 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_758
timestamp 1669390400
transform 1 0 86240 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_764
timestamp 1669390400
transform 1 0 86912 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_768
timestamp 1669390400
transform 1 0 87360 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_775
timestamp 1669390400
transform 1 0 88144 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_806
timestamp 1669390400
transform 1 0 91616 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_808
timestamp 1669390400
transform 1 0 91840 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_811
timestamp 1669390400
transform 1 0 92176 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_815
timestamp 1669390400
transform 1 0 92624 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_818
timestamp 1669390400
transform 1 0 92960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_70_821
timestamp 1669390400
transform 1 0 93296 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_829
timestamp 1669390400
transform 1 0 94192 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_831
timestamp 1669390400
transform 1 0 94416 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_837
timestamp 1669390400
transform 1 0 95088 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_844
timestamp 1669390400
transform 1 0 95872 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_851
timestamp 1669390400
transform 1 0 96656 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_855
timestamp 1669390400
transform 1 0 97104 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_859
timestamp 1669390400
transform 1 0 97552 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_863
timestamp 1669390400
transform 1 0 98000 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_865
timestamp 1669390400
transform 1 0 98224 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_66
timestamp 1669390400
transform 1 0 8736 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1669390400
transform 1 0 9184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1669390400
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_137
timestamp 1669390400
transform 1 0 16688 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1669390400
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1669390400
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_208
timestamp 1669390400
transform 1 0 24640 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1669390400
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1669390400
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_279
timestamp 1669390400
transform 1 0 32592 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1669390400
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1669390400
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_350
timestamp 1669390400
transform 1 0 40544 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_357
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_389
timestamp 1669390400
transform 1 0 44912 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_405
timestamp 1669390400
transform 1 0 46704 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_409
timestamp 1669390400
transform 1 0 47152 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_417
timestamp 1669390400
transform 1 0 48048 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1669390400
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_428
timestamp 1669390400
transform 1 0 49280 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_458
timestamp 1669390400
transform 1 0 52640 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_462
timestamp 1669390400
transform 1 0 53088 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_466
timestamp 1669390400
transform 1 0 53536 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1669390400
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_499
timestamp 1669390400
transform 1 0 57232 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_505
timestamp 1669390400
transform 1 0 57904 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_512
timestamp 1669390400
transform 1 0 58688 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_516
timestamp 1669390400
transform 1 0 59136 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_547
timestamp 1669390400
transform 1 0 62608 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_554
timestamp 1669390400
transform 1 0 63392 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_561
timestamp 1669390400
transform 1 0 64176 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_565
timestamp 1669390400
transform 1 0 64624 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_567
timestamp 1669390400
transform 1 0 64848 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_570
timestamp 1669390400
transform 1 0 65184 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_572
timestamp 1669390400
transform 1 0 65408 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_605
timestamp 1669390400
transform 1 0 69104 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_609
timestamp 1669390400
transform 1 0 69552 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_613
timestamp 1669390400
transform 1 0 70000 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_620
timestamp 1669390400
transform 1 0 70784 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_628
timestamp 1669390400
transform 1 0 71680 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1669390400
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_641
timestamp 1669390400
transform 1 0 73136 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_682
timestamp 1669390400
transform 1 0 77728 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_690
timestamp 1669390400
transform 1 0 78624 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_698
timestamp 1669390400
transform 1 0 79520 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_702
timestamp 1669390400
transform 1 0 79968 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_706
timestamp 1669390400
transform 1 0 80416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_712
timestamp 1669390400
transform 1 0 81088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_715
timestamp 1669390400
transform 1 0 81424 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_719
timestamp 1669390400
transform 1 0 81872 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_723
timestamp 1669390400
transform 1 0 82320 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_727
timestamp 1669390400
transform 1 0 82768 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_731
timestamp 1669390400
transform 1 0 83216 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_735
timestamp 1669390400
transform 1 0 83664 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_739
timestamp 1669390400
transform 1 0 84112 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_743
timestamp 1669390400
transform 1 0 84560 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_747
timestamp 1669390400
transform 1 0 85008 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_751
timestamp 1669390400
transform 1 0 85456 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_755
timestamp 1669390400
transform 1 0 85904 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_771
timestamp 1669390400
transform 1 0 87696 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_779
timestamp 1669390400
transform 1 0 88592 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_783
timestamp 1669390400
transform 1 0 89040 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_785
timestamp 1669390400
transform 1 0 89264 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_791
timestamp 1669390400
transform 1 0 89936 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_799
timestamp 1669390400
transform 1 0 90832 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_803
timestamp 1669390400
transform 1 0 91280 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_805
timestamp 1669390400
transform 1 0 91504 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_71_808
timestamp 1669390400
transform 1 0 91840 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_824
timestamp 1669390400
transform 1 0 93632 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_828
timestamp 1669390400
transform 1 0 94080 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_71_834
timestamp 1669390400
transform 1 0 94752 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_838
timestamp 1669390400
transform 1 0 95200 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_840
timestamp 1669390400
transform 1 0 95424 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_846
timestamp 1669390400
transform 1 0 96096 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_850
timestamp 1669390400
transform 1 0 96544 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_854
timestamp 1669390400
transform 1 0 96992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_857
timestamp 1669390400
transform 1 0 97328 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_865
timestamp 1669390400
transform 1 0 98224 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1669390400
transform 1 0 5152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1669390400
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_101
timestamp 1669390400
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1669390400
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1669390400
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_172
timestamp 1669390400
transform 1 0 20608 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1669390400
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1669390400
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_243
timestamp 1669390400
transform 1 0 28560 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1669390400
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1669390400
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_314
timestamp 1669390400
transform 1 0 36512 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1669390400
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1669390400
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_385
timestamp 1669390400
transform 1 0 44464 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1669390400
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_392
timestamp 1669390400
transform 1 0 45248 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_72_408
timestamp 1669390400
transform 1 0 47040 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_416
timestamp 1669390400
transform 1 0 47936 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_447
timestamp 1669390400
transform 1 0 51408 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_451
timestamp 1669390400
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_455
timestamp 1669390400
transform 1 0 52304 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_457
timestamp 1669390400
transform 1 0 52528 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1669390400
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_463
timestamp 1669390400
transform 1 0 53200 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_465
timestamp 1669390400
transform 1 0 53424 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_495
timestamp 1669390400
transform 1 0 56784 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_502
timestamp 1669390400
transform 1 0 57568 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_506
timestamp 1669390400
transform 1 0 58016 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_512
timestamp 1669390400
transform 1 0 58688 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_516
timestamp 1669390400
transform 1 0 59136 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_534
timestamp 1669390400
transform 1 0 61152 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_540
timestamp 1669390400
transform 1 0 61824 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_544
timestamp 1669390400
transform 1 0 62272 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_578
timestamp 1669390400
transform 1 0 66080 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_582
timestamp 1669390400
transform 1 0 66528 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_586
timestamp 1669390400
transform 1 0 66976 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_590
timestamp 1669390400
transform 1 0 67424 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_597
timestamp 1669390400
transform 1 0 68208 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_601
timestamp 1669390400
transform 1 0 68656 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_605
timestamp 1669390400
transform 1 0 69104 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_613
timestamp 1669390400
transform 1 0 70000 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_615
timestamp 1669390400
transform 1 0 70224 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_622
timestamp 1669390400
transform 1 0 71008 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_632
timestamp 1669390400
transform 1 0 72128 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_642
timestamp 1669390400
transform 1 0 73248 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_662
timestamp 1669390400
transform 1 0 75488 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_672
timestamp 1669390400
transform 1 0 76608 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_676
timestamp 1669390400
transform 1 0 77056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_683
timestamp 1669390400
transform 1 0 77840 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_691
timestamp 1669390400
transform 1 0 78736 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_695
timestamp 1669390400
transform 1 0 79184 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_728
timestamp 1669390400
transform 1 0 82880 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_732
timestamp 1669390400
transform 1 0 83328 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_736
timestamp 1669390400
transform 1 0 83776 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_740
timestamp 1669390400
transform 1 0 84224 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_744
timestamp 1669390400
transform 1 0 84672 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_747
timestamp 1669390400
transform 1 0 85008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_780
timestamp 1669390400
transform 1 0 88704 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_784
timestamp 1669390400
transform 1 0 89152 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_788
timestamp 1669390400
transform 1 0 89600 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_792
timestamp 1669390400
transform 1 0 90048 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_808
timestamp 1669390400
transform 1 0 91840 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_815
timestamp 1669390400
transform 1 0 92624 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_818
timestamp 1669390400
transform 1 0 92960 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_851
timestamp 1669390400
transform 1 0 96656 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_858
timestamp 1669390400
transform 1 0 97440 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_865
timestamp 1669390400
transform 1 0 98224 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_2
timestamp 1669390400
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_66
timestamp 1669390400
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_70
timestamp 1669390400
transform 1 0 9184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1669390400
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_137
timestamp 1669390400
transform 1 0 16688 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1669390400
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1669390400
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_208
timestamp 1669390400
transform 1 0 24640 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1669390400
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1669390400
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_279
timestamp 1669390400
transform 1 0 32592 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1669390400
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1669390400
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_350
timestamp 1669390400
transform 1 0 40544 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1669390400
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_357
timestamp 1669390400
transform 1 0 41328 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_389
timestamp 1669390400
transform 1 0 44912 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_405
timestamp 1669390400
transform 1 0 46704 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_413
timestamp 1669390400
transform 1 0 47600 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_417
timestamp 1669390400
transform 1 0 48048 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1669390400
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_428
timestamp 1669390400
transform 1 0 49280 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_445
timestamp 1669390400
transform 1 0 51184 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_449
timestamp 1669390400
transform 1 0 51632 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_453
timestamp 1669390400
transform 1 0 52080 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_469
timestamp 1669390400
transform 1 0 53872 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_477
timestamp 1669390400
transform 1 0 54768 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_486
timestamp 1669390400
transform 1 0 55776 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_493
timestamp 1669390400
transform 1 0 56560 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_499
timestamp 1669390400
transform 1 0 57232 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_502
timestamp 1669390400
transform 1 0 57568 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_73_506
timestamp 1669390400
transform 1 0 58016 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_522
timestamp 1669390400
transform 1 0 59808 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_530
timestamp 1669390400
transform 1 0 60704 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_534
timestamp 1669390400
transform 1 0 61152 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1669390400
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_570
timestamp 1669390400
transform 1 0 65184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_573
timestamp 1669390400
transform 1 0 65520 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_577
timestamp 1669390400
transform 1 0 65968 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_581
timestamp 1669390400
transform 1 0 66416 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_585
timestamp 1669390400
transform 1 0 66864 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_593
timestamp 1669390400
transform 1 0 67760 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_595
timestamp 1669390400
transform 1 0 67984 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_602
timestamp 1669390400
transform 1 0 68768 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_609
timestamp 1669390400
transform 1 0 69552 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_619
timestamp 1669390400
transform 1 0 70672 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_627
timestamp 1669390400
transform 1 0 71568 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_629
timestamp 1669390400
transform 1 0 71792 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_638
timestamp 1669390400
transform 1 0 72800 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_641
timestamp 1669390400
transform 1 0 73136 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_693
timestamp 1669390400
transform 1 0 78960 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_701
timestamp 1669390400
transform 1 0 79856 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_709
timestamp 1669390400
transform 1 0 80752 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_712
timestamp 1669390400
transform 1 0 81088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_717
timestamp 1669390400
transform 1 0 81648 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_721
timestamp 1669390400
transform 1 0 82096 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_725
timestamp 1669390400
transform 1 0 82544 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_729
timestamp 1669390400
transform 1 0 82992 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_733
timestamp 1669390400
transform 1 0 83440 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_742
timestamp 1669390400
transform 1 0 84448 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_776
timestamp 1669390400
transform 1 0 88256 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_780
timestamp 1669390400
transform 1 0 88704 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_783
timestamp 1669390400
transform 1 0 89040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_786
timestamp 1669390400
transform 1 0 89376 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_790
timestamp 1669390400
transform 1 0 89824 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_794
timestamp 1669390400
transform 1 0 90272 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_796
timestamp 1669390400
transform 1 0 90496 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_799
timestamp 1669390400
transform 1 0 90832 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_851
timestamp 1669390400
transform 1 0 96656 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_854
timestamp 1669390400
transform 1 0 96992 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_73_862
timestamp 1669390400
transform 1 0 97888 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_2
timestamp 1669390400
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_34
timestamp 1669390400
transform 1 0 5152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1669390400
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_101
timestamp 1669390400
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1669390400
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1669390400
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_172
timestamp 1669390400
transform 1 0 20608 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1669390400
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1669390400
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_243
timestamp 1669390400
transform 1 0 28560 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1669390400
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1669390400
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_314
timestamp 1669390400
transform 1 0 36512 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1669390400
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1669390400
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_385
timestamp 1669390400
transform 1 0 44464 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1669390400
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_392
timestamp 1669390400
transform 1 0 45248 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_408
timestamp 1669390400
transform 1 0 47040 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_416
timestamp 1669390400
transform 1 0 47936 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_420
timestamp 1669390400
transform 1 0 48384 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_422
timestamp 1669390400
transform 1 0 48608 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_425
timestamp 1669390400
transform 1 0 48944 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_442
timestamp 1669390400
transform 1 0 50848 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_446
timestamp 1669390400
transform 1 0 51296 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_454
timestamp 1669390400
transform 1 0 52192 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_458
timestamp 1669390400
transform 1 0 52640 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1669390400
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_463
timestamp 1669390400
transform 1 0 53200 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_466
timestamp 1669390400
transform 1 0 53536 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_474
timestamp 1669390400
transform 1 0 54432 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_483
timestamp 1669390400
transform 1 0 55440 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_487
timestamp 1669390400
transform 1 0 55888 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_491
timestamp 1669390400
transform 1 0 56336 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_507
timestamp 1669390400
transform 1 0 58128 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_509
timestamp 1669390400
transform 1 0 58352 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_512
timestamp 1669390400
transform 1 0 58688 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_519
timestamp 1669390400
transform 1 0 59472 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_523
timestamp 1669390400
transform 1 0 59920 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_527
timestamp 1669390400
transform 1 0 60368 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1669390400
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_534
timestamp 1669390400
transform 1 0 61152 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_538
timestamp 1669390400
transform 1 0 61600 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_571
timestamp 1669390400
transform 1 0 65296 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_575
timestamp 1669390400
transform 1 0 65744 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_579
timestamp 1669390400
transform 1 0 66192 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_587
timestamp 1669390400
transform 1 0 67088 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_597
timestamp 1669390400
transform 1 0 68208 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_601
timestamp 1669390400
transform 1 0 68656 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_605
timestamp 1669390400
transform 1 0 69104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_608
timestamp 1669390400
transform 1 0 69440 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_619
timestamp 1669390400
transform 1 0 70672 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_629
timestamp 1669390400
transform 1 0 71792 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_640
timestamp 1669390400
transform 1 0 73024 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_656
timestamp 1669390400
transform 1 0 74816 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_667
timestamp 1669390400
transform 1 0 76048 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_671
timestamp 1669390400
transform 1 0 76496 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1669390400
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_676
timestamp 1669390400
transform 1 0 77056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_685
timestamp 1669390400
transform 1 0 78064 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_695
timestamp 1669390400
transform 1 0 79184 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_702
timestamp 1669390400
transform 1 0 79968 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_712
timestamp 1669390400
transform 1 0 81088 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_720
timestamp 1669390400
transform 1 0 81984 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_724
timestamp 1669390400
transform 1 0 82432 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_728
timestamp 1669390400
transform 1 0 82880 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_730
timestamp 1669390400
transform 1 0 83104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_739
timestamp 1669390400
transform 1 0 84112 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_743
timestamp 1669390400
transform 1 0 84560 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_747
timestamp 1669390400
transform 1 0 85008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_756
timestamp 1669390400
transform 1 0 86016 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_760
timestamp 1669390400
transform 1 0 86464 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_764
timestamp 1669390400
transform 1 0 86912 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_768
timestamp 1669390400
transform 1 0 87360 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_772
timestamp 1669390400
transform 1 0 87808 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_782
timestamp 1669390400
transform 1 0 88928 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_786
timestamp 1669390400
transform 1 0 89376 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_790
timestamp 1669390400
transform 1 0 89824 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_806
timestamp 1669390400
transform 1 0 91616 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_814
timestamp 1669390400
transform 1 0 92512 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_818
timestamp 1669390400
transform 1 0 92960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_821
timestamp 1669390400
transform 1 0 93296 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_74_854
timestamp 1669390400
transform 1 0 96992 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_862
timestamp 1669390400
transform 1 0 97888 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_2
timestamp 1669390400
transform 1 0 1568 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_5
timestamp 1669390400
transform 1 0 1904 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_69
timestamp 1669390400
transform 1 0 9072 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1669390400
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_137
timestamp 1669390400
transform 1 0 16688 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1669390400
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1669390400
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_208
timestamp 1669390400
transform 1 0 24640 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1669390400
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1669390400
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_279
timestamp 1669390400
transform 1 0 32592 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1669390400
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1669390400
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_350
timestamp 1669390400
transform 1 0 40544 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1669390400
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_357
timestamp 1669390400
transform 1 0 41328 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_75_389
timestamp 1669390400
transform 1 0 44912 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_405
timestamp 1669390400
transform 1 0 46704 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_413
timestamp 1669390400
transform 1 0 47600 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_417
timestamp 1669390400
transform 1 0 48048 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1669390400
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_428
timestamp 1669390400
transform 1 0 49280 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_432
timestamp 1669390400
transform 1 0 49728 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_484
timestamp 1669390400
transform 1 0 55552 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_488
timestamp 1669390400
transform 1 0 56000 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_492
timestamp 1669390400
transform 1 0 56448 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1669390400
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_499
timestamp 1669390400
transform 1 0 57232 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_508
timestamp 1669390400
transform 1 0 58240 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_512
timestamp 1669390400
transform 1 0 58688 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_514
timestamp 1669390400
transform 1 0 58912 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_520
timestamp 1669390400
transform 1 0 59584 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_524
timestamp 1669390400
transform 1 0 60032 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_528
timestamp 1669390400
transform 1 0 60480 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_536
timestamp 1669390400
transform 1 0 61376 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_538
timestamp 1669390400
transform 1 0 61600 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_547
timestamp 1669390400
transform 1 0 62608 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_557
timestamp 1669390400
transform 1 0 63728 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_561
timestamp 1669390400
transform 1 0 64176 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_565
timestamp 1669390400
transform 1 0 64624 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1669390400
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_570
timestamp 1669390400
transform 1 0 65184 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_574
timestamp 1669390400
transform 1 0 65632 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_577
timestamp 1669390400
transform 1 0 65968 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_608
timestamp 1669390400
transform 1 0 69440 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_616
timestamp 1669390400
transform 1 0 70336 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_628
timestamp 1669390400
transform 1 0 71680 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1669390400
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_641
timestamp 1669390400
transform 1 0 73136 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_682
timestamp 1669390400
transform 1 0 77728 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_690
timestamp 1669390400
transform 1 0 78624 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_694
timestamp 1669390400
transform 1 0 79072 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_702
timestamp 1669390400
transform 1 0 79968 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_706
timestamp 1669390400
transform 1 0 80416 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_712
timestamp 1669390400
transform 1 0 81088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_721
timestamp 1669390400
transform 1 0 82096 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_729
timestamp 1669390400
transform 1 0 82992 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_733
timestamp 1669390400
transform 1 0 83440 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_737
timestamp 1669390400
transform 1 0 83888 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_746
timestamp 1669390400
transform 1 0 84896 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_750
timestamp 1669390400
transform 1 0 85344 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_754
timestamp 1669390400
transform 1 0 85792 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_764
timestamp 1669390400
transform 1 0 86912 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_774
timestamp 1669390400
transform 1 0 88032 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_778
timestamp 1669390400
transform 1 0 88480 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_780
timestamp 1669390400
transform 1 0 88704 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_783
timestamp 1669390400
transform 1 0 89040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_816
timestamp 1669390400
transform 1 0 92736 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_820
timestamp 1669390400
transform 1 0 93184 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_851
timestamp 1669390400
transform 1 0 96656 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_854
timestamp 1669390400
transform 1 0 96992 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_75_862
timestamp 1669390400
transform 1 0 97888 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_2
timestamp 1669390400
transform 1 0 1568 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_9
timestamp 1669390400
transform 1 0 2352 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_76_25
timestamp 1669390400
transform 1 0 4144 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_33
timestamp 1669390400
transform 1 0 5040 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1669390400
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_101
timestamp 1669390400
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1669390400
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1669390400
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_172
timestamp 1669390400
transform 1 0 20608 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1669390400
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1669390400
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_243
timestamp 1669390400
transform 1 0 28560 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1669390400
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1669390400
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_314
timestamp 1669390400
transform 1 0 36512 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1669390400
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1669390400
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_385
timestamp 1669390400
transform 1 0 44464 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1669390400
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_392
timestamp 1669390400
transform 1 0 45248 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_424
timestamp 1669390400
transform 1 0 48832 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_426
timestamp 1669390400
transform 1 0 49056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_456
timestamp 1669390400
transform 1 0 52416 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1669390400
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_463
timestamp 1669390400
transform 1 0 53200 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_465
timestamp 1669390400
transform 1 0 53424 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_498
timestamp 1669390400
transform 1 0 57120 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_502
timestamp 1669390400
transform 1 0 57568 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_515
timestamp 1669390400
transform 1 0 59024 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_526
timestamp 1669390400
transform 1 0 60256 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_530
timestamp 1669390400
transform 1 0 60704 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_534
timestamp 1669390400
transform 1 0 61152 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_538
timestamp 1669390400
transform 1 0 61600 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_548
timestamp 1669390400
transform 1 0 62720 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_552
timestamp 1669390400
transform 1 0 63168 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_556
timestamp 1669390400
transform 1 0 63616 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_572
timestamp 1669390400
transform 1 0 65408 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_574
timestamp 1669390400
transform 1 0 65632 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_577
timestamp 1669390400
transform 1 0 65968 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_581
timestamp 1669390400
transform 1 0 66416 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_585
timestamp 1669390400
transform 1 0 66864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_592
timestamp 1669390400
transform 1 0 67648 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1669390400
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_605
timestamp 1669390400
transform 1 0 69104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_608
timestamp 1669390400
transform 1 0 69440 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_616
timestamp 1669390400
transform 1 0 70336 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_620
timestamp 1669390400
transform 1 0 70784 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_624
timestamp 1669390400
transform 1 0 71232 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_634
timestamp 1669390400
transform 1 0 72352 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1669390400
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_676
timestamp 1669390400
transform 1 0 77056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_685
timestamp 1669390400
transform 1 0 78064 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_693
timestamp 1669390400
transform 1 0 78960 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_727
timestamp 1669390400
transform 1 0 82768 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_731
timestamp 1669390400
transform 1 0 83216 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_741
timestamp 1669390400
transform 1 0 84336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_747
timestamp 1669390400
transform 1 0 85008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_750
timestamp 1669390400
transform 1 0 85344 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_752
timestamp 1669390400
transform 1 0 85568 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_762
timestamp 1669390400
transform 1 0 86688 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_766
timestamp 1669390400
transform 1 0 87136 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_770
timestamp 1669390400
transform 1 0 87584 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_772
timestamp 1669390400
transform 1 0 87808 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_805
timestamp 1669390400
transform 1 0 91504 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_809
timestamp 1669390400
transform 1 0 91952 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_813
timestamp 1669390400
transform 1 0 92400 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_815
timestamp 1669390400
transform 1 0 92624 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_818
timestamp 1669390400
transform 1 0 92960 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_822
timestamp 1669390400
transform 1 0 93408 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_825
timestamp 1669390400
transform 1 0 93744 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_832
timestamp 1669390400
transform 1 0 94528 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_839
timestamp 1669390400
transform 1 0 95312 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_843
timestamp 1669390400
transform 1 0 95760 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_847
timestamp 1669390400
transform 1 0 96208 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_863
timestamp 1669390400
transform 1 0 98000 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_865
timestamp 1669390400
transform 1 0 98224 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_2
timestamp 1669390400
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_66
timestamp 1669390400
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_70
timestamp 1669390400
transform 1 0 9184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1669390400
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_137
timestamp 1669390400
transform 1 0 16688 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1669390400
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1669390400
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_208
timestamp 1669390400
transform 1 0 24640 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1669390400
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1669390400
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_279
timestamp 1669390400
transform 1 0 32592 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1669390400
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1669390400
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_350
timestamp 1669390400
transform 1 0 40544 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1669390400
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1669390400
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_421
timestamp 1669390400
transform 1 0 48496 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1669390400
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_428
timestamp 1669390400
transform 1 0 49280 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_458
timestamp 1669390400
transform 1 0 52640 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_462
timestamp 1669390400
transform 1 0 53088 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1669390400
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_499
timestamp 1669390400
transform 1 0 57232 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_532
timestamp 1669390400
transform 1 0 60928 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_536
timestamp 1669390400
transform 1 0 61376 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_77_540
timestamp 1669390400
transform 1 0 61824 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_556
timestamp 1669390400
transform 1 0 63616 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_564
timestamp 1669390400
transform 1 0 64512 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_570
timestamp 1669390400
transform 1 0 65184 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_580
timestamp 1669390400
transform 1 0 66304 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_614
timestamp 1669390400
transform 1 0 70112 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_616
timestamp 1669390400
transform 1 0 70336 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_623
timestamp 1669390400
transform 1 0 71120 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_627
timestamp 1669390400
transform 1 0 71568 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1669390400
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_641
timestamp 1669390400
transform 1 0 73136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_679
timestamp 1669390400
transform 1 0 77392 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_690
timestamp 1669390400
transform 1 0 78624 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_698
timestamp 1669390400
transform 1 0 79520 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_706
timestamp 1669390400
transform 1 0 80416 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_712
timestamp 1669390400
transform 1 0 81088 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_714
timestamp 1669390400
transform 1 0 81312 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_724
timestamp 1669390400
transform 1 0 82432 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_735
timestamp 1669390400
transform 1 0 83664 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_739
timestamp 1669390400
transform 1 0 84112 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_743
timestamp 1669390400
transform 1 0 84560 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_750
timestamp 1669390400
transform 1 0 85344 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_754
timestamp 1669390400
transform 1 0 85792 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_763
timestamp 1669390400
transform 1 0 86800 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_767
timestamp 1669390400
transform 1 0 87248 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_771
timestamp 1669390400
transform 1 0 87696 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_775
timestamp 1669390400
transform 1 0 88144 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_779
timestamp 1669390400
transform 1 0 88592 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_783
timestamp 1669390400
transform 1 0 89040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_816
timestamp 1669390400
transform 1 0 92736 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_820
timestamp 1669390400
transform 1 0 93184 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_824
timestamp 1669390400
transform 1 0 93632 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_834
timestamp 1669390400
transform 1 0 94752 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_851
timestamp 1669390400
transform 1 0 96656 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_854
timestamp 1669390400
transform 1 0 96992 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_77_862
timestamp 1669390400
transform 1 0 97888 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_2
timestamp 1669390400
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_34
timestamp 1669390400
transform 1 0 5152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1669390400
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_101
timestamp 1669390400
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1669390400
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1669390400
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_172
timestamp 1669390400
transform 1 0 20608 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1669390400
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1669390400
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_243
timestamp 1669390400
transform 1 0 28560 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1669390400
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1669390400
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_314
timestamp 1669390400
transform 1 0 36512 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1669390400
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1669390400
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_385
timestamp 1669390400
transform 1 0 44464 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1669390400
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_392
timestamp 1669390400
transform 1 0 45248 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_408
timestamp 1669390400
transform 1 0 47040 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_416
timestamp 1669390400
transform 1 0 47936 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_420
timestamp 1669390400
transform 1 0 48384 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_451
timestamp 1669390400
transform 1 0 51856 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_458
timestamp 1669390400
transform 1 0 52640 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1669390400
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_463
timestamp 1669390400
transform 1 0 53200 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_469
timestamp 1669390400
transform 1 0 53872 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_473
timestamp 1669390400
transform 1 0 54320 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_477
timestamp 1669390400
transform 1 0 54768 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_481
timestamp 1669390400
transform 1 0 55216 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_485
timestamp 1669390400
transform 1 0 55664 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_498
timestamp 1669390400
transform 1 0 57120 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_508
timestamp 1669390400
transform 1 0 58240 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_512
timestamp 1669390400
transform 1 0 58688 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_516
timestamp 1669390400
transform 1 0 59136 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_520
timestamp 1669390400
transform 1 0 59584 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_524
timestamp 1669390400
transform 1 0 60032 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1669390400
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_534
timestamp 1669390400
transform 1 0 61152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_537
timestamp 1669390400
transform 1 0 61488 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_541
timestamp 1669390400
transform 1 0 61936 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_557
timestamp 1669390400
transform 1 0 63728 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_587
timestamp 1669390400
transform 1 0 67088 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_591
timestamp 1669390400
transform 1 0 67536 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_594
timestamp 1669390400
transform 1 0 67872 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_598
timestamp 1669390400
transform 1 0 68320 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_602
timestamp 1669390400
transform 1 0 68768 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_605
timestamp 1669390400
transform 1 0 69104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_612
timestamp 1669390400
transform 1 0 69888 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_622
timestamp 1669390400
transform 1 0 71008 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_629
timestamp 1669390400
transform 1 0 71792 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_633
timestamp 1669390400
transform 1 0 72240 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_635
timestamp 1669390400
transform 1 0 72464 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_673
timestamp 1669390400
transform 1 0 76720 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_676
timestamp 1669390400
transform 1 0 77056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_679
timestamp 1669390400
transform 1 0 77392 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_681
timestamp 1669390400
transform 1 0 77616 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_688
timestamp 1669390400
transform 1 0 78400 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_698
timestamp 1669390400
transform 1 0 79520 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_706
timestamp 1669390400
transform 1 0 80416 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_713
timestamp 1669390400
transform 1 0 81200 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_717
timestamp 1669390400
transform 1 0 81648 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_721
timestamp 1669390400
transform 1 0 82096 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_725
timestamp 1669390400
transform 1 0 82544 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_729
timestamp 1669390400
transform 1 0 82992 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_733
timestamp 1669390400
transform 1 0 83440 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_742
timestamp 1669390400
transform 1 0 84448 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_744
timestamp 1669390400
transform 1 0 84672 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_747
timestamp 1669390400
transform 1 0 85008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_753
timestamp 1669390400
transform 1 0 85680 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_763
timestamp 1669390400
transform 1 0 86800 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_767
timestamp 1669390400
transform 1 0 87248 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_800
timestamp 1669390400
transform 1 0 90944 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_78_804
timestamp 1669390400
transform 1 0 91392 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_812
timestamp 1669390400
transform 1 0 92288 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_818
timestamp 1669390400
transform 1 0 92960 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_822
timestamp 1669390400
transform 1 0 93408 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_826
timestamp 1669390400
transform 1 0 93856 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_857
timestamp 1669390400
transform 1 0 97328 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_861
timestamp 1669390400
transform 1 0 97776 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_865
timestamp 1669390400
transform 1 0 98224 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_2
timestamp 1669390400
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_66
timestamp 1669390400
transform 1 0 8736 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_70
timestamp 1669390400
transform 1 0 9184 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1669390400
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_137
timestamp 1669390400
transform 1 0 16688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1669390400
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1669390400
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_208
timestamp 1669390400
transform 1 0 24640 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1669390400
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1669390400
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_279
timestamp 1669390400
transform 1 0 32592 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1669390400
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1669390400
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_350
timestamp 1669390400
transform 1 0 40544 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1669390400
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1669390400
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_421
timestamp 1669390400
transform 1 0 48496 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1669390400
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_428
timestamp 1669390400
transform 1 0 49280 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_458
timestamp 1669390400
transform 1 0 52640 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_465
timestamp 1669390400
transform 1 0 53424 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_467
timestamp 1669390400
transform 1 0 53648 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_473
timestamp 1669390400
transform 1 0 54320 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_477
timestamp 1669390400
transform 1 0 54768 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_484
timestamp 1669390400
transform 1 0 55552 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_488
timestamp 1669390400
transform 1 0 56000 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_492
timestamp 1669390400
transform 1 0 56448 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1669390400
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_499
timestamp 1669390400
transform 1 0 57232 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_508
timestamp 1669390400
transform 1 0 58240 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_515
timestamp 1669390400
transform 1 0 59024 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_519
timestamp 1669390400
transform 1 0 59472 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_521
timestamp 1669390400
transform 1 0 59696 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_551
timestamp 1669390400
transform 1 0 63056 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_555
timestamp 1669390400
transform 1 0 63504 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_559
timestamp 1669390400
transform 1 0 63952 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1669390400
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_570
timestamp 1669390400
transform 1 0 65184 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_621
timestamp 1669390400
transform 1 0 70896 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_625
timestamp 1669390400
transform 1 0 71344 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_629
timestamp 1669390400
transform 1 0 71792 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_633
timestamp 1669390400
transform 1 0 72240 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_635
timestamp 1669390400
transform 1 0 72464 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_638
timestamp 1669390400
transform 1 0 72800 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_641
timestamp 1669390400
transform 1 0 73136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_679
timestamp 1669390400
transform 1 0 77392 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_687
timestamp 1669390400
transform 1 0 78288 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_689
timestamp 1669390400
transform 1 0 78512 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_696
timestamp 1669390400
transform 1 0 79296 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_703
timestamp 1669390400
transform 1 0 80080 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_707
timestamp 1669390400
transform 1 0 80528 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_709
timestamp 1669390400
transform 1 0 80752 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_712
timestamp 1669390400
transform 1 0 81088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_715
timestamp 1669390400
transform 1 0 81424 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_719
timestamp 1669390400
transform 1 0 81872 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_723
timestamp 1669390400
transform 1 0 82320 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_727
timestamp 1669390400
transform 1 0 82768 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_758
timestamp 1669390400
transform 1 0 86240 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_765
timestamp 1669390400
transform 1 0 87024 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_769
timestamp 1669390400
transform 1 0 87472 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_771
timestamp 1669390400
transform 1 0 87696 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_777
timestamp 1669390400
transform 1 0 88368 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_783
timestamp 1669390400
transform 1 0 89040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_789
timestamp 1669390400
transform 1 0 89712 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_796
timestamp 1669390400
transform 1 0 90496 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_800
timestamp 1669390400
transform 1 0 90944 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_79_804
timestamp 1669390400
transform 1 0 91392 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_820
timestamp 1669390400
transform 1 0 93184 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_826
timestamp 1669390400
transform 1 0 93856 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_834
timestamp 1669390400
transform 1 0 94752 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_851
timestamp 1669390400
transform 1 0 96656 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_854
timestamp 1669390400
transform 1 0 96992 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_79_862
timestamp 1669390400
transform 1 0 97888 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_2
timestamp 1669390400
transform 1 0 1568 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_34
timestamp 1669390400
transform 1 0 5152 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1669390400
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_101
timestamp 1669390400
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1669390400
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1669390400
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_172
timestamp 1669390400
transform 1 0 20608 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1669390400
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1669390400
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_243
timestamp 1669390400
transform 1 0 28560 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1669390400
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1669390400
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_314
timestamp 1669390400
transform 1 0 36512 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1669390400
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1669390400
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_385
timestamp 1669390400
transform 1 0 44464 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1669390400
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_392
timestamp 1669390400
transform 1 0 45248 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_424
timestamp 1669390400
transform 1 0 48832 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_431
timestamp 1669390400
transform 1 0 49616 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_438
timestamp 1669390400
transform 1 0 50400 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_445
timestamp 1669390400
transform 1 0 51184 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_452
timestamp 1669390400
transform 1 0 51968 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_459
timestamp 1669390400
transform 1 0 52752 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_463
timestamp 1669390400
transform 1 0 53200 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_494
timestamp 1669390400
transform 1 0 56672 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_498
timestamp 1669390400
transform 1 0 57120 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_506
timestamp 1669390400
transform 1 0 58016 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_509
timestamp 1669390400
transform 1 0 58352 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_516
timestamp 1669390400
transform 1 0 59136 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_520
timestamp 1669390400
transform 1 0 59584 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_524
timestamp 1669390400
transform 1 0 60032 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1669390400
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_534
timestamp 1669390400
transform 1 0 61152 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_551
timestamp 1669390400
transform 1 0 63056 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_80_555
timestamp 1669390400
transform 1 0 63504 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_563
timestamp 1669390400
transform 1 0 64400 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_567
timestamp 1669390400
transform 1 0 64848 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_570
timestamp 1669390400
transform 1 0 65184 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_587
timestamp 1669390400
transform 1 0 67088 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_598
timestamp 1669390400
transform 1 0 68320 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1669390400
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_605
timestamp 1669390400
transform 1 0 69104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_611
timestamp 1669390400
transform 1 0 69776 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_615
timestamp 1669390400
transform 1 0 70224 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_618
timestamp 1669390400
transform 1 0 70560 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_622
timestamp 1669390400
transform 1 0 71008 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_626
timestamp 1669390400
transform 1 0 71456 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_630
timestamp 1669390400
transform 1 0 71904 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_634
timestamp 1669390400
transform 1 0 72352 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_643
timestamp 1669390400
transform 1 0 73360 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_651
timestamp 1669390400
transform 1 0 74256 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_659
timestamp 1669390400
transform 1 0 75152 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_667
timestamp 1669390400
transform 1 0 76048 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_671
timestamp 1669390400
transform 1 0 76496 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1669390400
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_676
timestamp 1669390400
transform 1 0 77056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_683
timestamp 1669390400
transform 1 0 77840 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_687
timestamp 1669390400
transform 1 0 78288 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_717
timestamp 1669390400
transform 1 0 81648 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_721
timestamp 1669390400
transform 1 0 82096 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_725
timestamp 1669390400
transform 1 0 82544 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_729
timestamp 1669390400
transform 1 0 82992 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_733
timestamp 1669390400
transform 1 0 83440 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_736
timestamp 1669390400
transform 1 0 83776 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_743
timestamp 1669390400
transform 1 0 84560 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_747
timestamp 1669390400
transform 1 0 85008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_750
timestamp 1669390400
transform 1 0 85344 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_752
timestamp 1669390400
transform 1 0 85568 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_758
timestamp 1669390400
transform 1 0 86240 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_762
timestamp 1669390400
transform 1 0 86688 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_795
timestamp 1669390400
transform 1 0 90384 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_802
timestamp 1669390400
transform 1 0 91168 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_806
timestamp 1669390400
transform 1 0 91616 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_810
timestamp 1669390400
transform 1 0 92064 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_812
timestamp 1669390400
transform 1 0 92288 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_815
timestamp 1669390400
transform 1 0 92624 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_818
timestamp 1669390400
transform 1 0 92960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_825
timestamp 1669390400
transform 1 0 93744 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_827
timestamp 1669390400
transform 1 0 93968 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_830
timestamp 1669390400
transform 1 0 94304 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_861
timestamp 1669390400
transform 1 0 97776 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_865
timestamp 1669390400
transform 1 0 98224 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_2
timestamp 1669390400
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_66
timestamp 1669390400
transform 1 0 8736 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_70
timestamp 1669390400
transform 1 0 9184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1669390400
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_137
timestamp 1669390400
transform 1 0 16688 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1669390400
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1669390400
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_208
timestamp 1669390400
transform 1 0 24640 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1669390400
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1669390400
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_279
timestamp 1669390400
transform 1 0 32592 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1669390400
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1669390400
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_350
timestamp 1669390400
transform 1 0 40544 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1669390400
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_357
timestamp 1669390400
transform 1 0 41328 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_389
timestamp 1669390400
transform 1 0 44912 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_405
timestamp 1669390400
transform 1 0 46704 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_413
timestamp 1669390400
transform 1 0 47600 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_417
timestamp 1669390400
transform 1 0 48048 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_421
timestamp 1669390400
transform 1 0 48496 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1669390400
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_428
timestamp 1669390400
transform 1 0 49280 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_430
timestamp 1669390400
transform 1 0 49504 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_433
timestamp 1669390400
transform 1 0 49840 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_440
timestamp 1669390400
transform 1 0 50624 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_442
timestamp 1669390400
transform 1 0 50848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_448
timestamp 1669390400
transform 1 0 51520 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_455
timestamp 1669390400
transform 1 0 52304 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_462
timestamp 1669390400
transform 1 0 53088 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_466
timestamp 1669390400
transform 1 0 53536 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_470
timestamp 1669390400
transform 1 0 53984 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_81_474
timestamp 1669390400
transform 1 0 54432 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_490
timestamp 1669390400
transform 1 0 56224 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_494
timestamp 1669390400
transform 1 0 56672 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1669390400
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_499
timestamp 1669390400
transform 1 0 57232 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_507
timestamp 1669390400
transform 1 0 58128 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_513
timestamp 1669390400
transform 1 0 58800 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_517
timestamp 1669390400
transform 1 0 59248 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_519
timestamp 1669390400
transform 1 0 59472 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_549
timestamp 1669390400
transform 1 0 62832 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_553
timestamp 1669390400
transform 1 0 63280 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_557
timestamp 1669390400
transform 1 0 63728 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_565
timestamp 1669390400
transform 1 0 64624 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1669390400
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_570
timestamp 1669390400
transform 1 0 65184 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_578
timestamp 1669390400
transform 1 0 66080 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_580
timestamp 1669390400
transform 1 0 66304 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_610
timestamp 1669390400
transform 1 0 69664 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_617
timestamp 1669390400
transform 1 0 70448 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_621
timestamp 1669390400
transform 1 0 70896 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_625
timestamp 1669390400
transform 1 0 71344 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_627
timestamp 1669390400
transform 1 0 71568 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_634
timestamp 1669390400
transform 1 0 72352 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1669390400
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_641
timestamp 1669390400
transform 1 0 73136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_650
timestamp 1669390400
transform 1 0 74144 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_658
timestamp 1669390400
transform 1 0 75040 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_662
timestamp 1669390400
transform 1 0 75488 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_664
timestamp 1669390400
transform 1 0 75712 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_670
timestamp 1669390400
transform 1 0 76384 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_678
timestamp 1669390400
transform 1 0 77280 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_709
timestamp 1669390400
transform 1 0 80752 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_712
timestamp 1669390400
transform 1 0 81088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_718
timestamp 1669390400
transform 1 0 81760 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_722
timestamp 1669390400
transform 1 0 82208 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_726
timestamp 1669390400
transform 1 0 82656 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_728
timestamp 1669390400
transform 1 0 82880 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_734
timestamp 1669390400
transform 1 0 83552 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_738
timestamp 1669390400
transform 1 0 84000 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_742
timestamp 1669390400
transform 1 0 84448 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_746
timestamp 1669390400
transform 1 0 84896 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_753
timestamp 1669390400
transform 1 0 85680 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_757
timestamp 1669390400
transform 1 0 86128 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_763
timestamp 1669390400
transform 1 0 86800 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_767
timestamp 1669390400
transform 1 0 87248 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_774
timestamp 1669390400
transform 1 0 88032 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_778
timestamp 1669390400
transform 1 0 88480 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_780
timestamp 1669390400
transform 1 0 88704 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_783
timestamp 1669390400
transform 1 0 89040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_834
timestamp 1669390400
transform 1 0 94752 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_851
timestamp 1669390400
transform 1 0 96656 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_854
timestamp 1669390400
transform 1 0 96992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_857
timestamp 1669390400
transform 1 0 97328 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_81_861
timestamp 1669390400
transform 1 0 97776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_865
timestamp 1669390400
transform 1 0 98224 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_2
timestamp 1669390400
transform 1 0 1568 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_34
timestamp 1669390400
transform 1 0 5152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1669390400
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_101
timestamp 1669390400
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1669390400
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1669390400
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_172
timestamp 1669390400
transform 1 0 20608 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1669390400
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1669390400
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_243
timestamp 1669390400
transform 1 0 28560 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1669390400
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1669390400
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_314
timestamp 1669390400
transform 1 0 36512 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1669390400
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1669390400
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_385
timestamp 1669390400
transform 1 0 44464 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1669390400
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_392
timestamp 1669390400
transform 1 0 45248 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_82_408
timestamp 1669390400
transform 1 0 47040 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_416
timestamp 1669390400
transform 1 0 47936 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_420
timestamp 1669390400
transform 1 0 48384 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_422
timestamp 1669390400
transform 1 0 48608 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_452
timestamp 1669390400
transform 1 0 51968 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_456
timestamp 1669390400
transform 1 0 52416 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1669390400
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_463
timestamp 1669390400
transform 1 0 53200 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_466
timestamp 1669390400
transform 1 0 53536 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_470
timestamp 1669390400
transform 1 0 53984 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_474
timestamp 1669390400
transform 1 0 54432 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_476
timestamp 1669390400
transform 1 0 54656 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_479
timestamp 1669390400
transform 1 0 54992 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_511
timestamp 1669390400
transform 1 0 58576 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_515
timestamp 1669390400
transform 1 0 59024 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_517
timestamp 1669390400
transform 1 0 59248 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_520
timestamp 1669390400
transform 1 0 59584 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_524
timestamp 1669390400
transform 1 0 60032 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1669390400
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_534
timestamp 1669390400
transform 1 0 61152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_550
timestamp 1669390400
transform 1 0 62944 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_554
timestamp 1669390400
transform 1 0 63392 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_558
timestamp 1669390400
transform 1 0 63840 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_588
timestamp 1669390400
transform 1 0 67200 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_595
timestamp 1669390400
transform 1 0 67984 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1669390400
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_605
timestamp 1669390400
transform 1 0 69104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_608
timestamp 1669390400
transform 1 0 69440 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_610
timestamp 1669390400
transform 1 0 69664 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_613
timestamp 1669390400
transform 1 0 70000 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_617
timestamp 1669390400
transform 1 0 70448 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_620
timestamp 1669390400
transform 1 0 70784 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_624
timestamp 1669390400
transform 1 0 71232 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_628
timestamp 1669390400
transform 1 0 71680 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_632
timestamp 1669390400
transform 1 0 72128 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_640
timestamp 1669390400
transform 1 0 73024 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_650
timestamp 1669390400
transform 1 0 74144 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_654
timestamp 1669390400
transform 1 0 74592 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_658
timestamp 1669390400
transform 1 0 75040 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_662
timestamp 1669390400
transform 1 0 75488 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_666
timestamp 1669390400
transform 1 0 75936 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_670
timestamp 1669390400
transform 1 0 76384 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_676
timestamp 1669390400
transform 1 0 77056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_727
timestamp 1669390400
transform 1 0 82768 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_731
timestamp 1669390400
transform 1 0 83216 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_738
timestamp 1669390400
transform 1 0 84000 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_742
timestamp 1669390400
transform 1 0 84448 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_744
timestamp 1669390400
transform 1 0 84672 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_747
timestamp 1669390400
transform 1 0 85008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_777
timestamp 1669390400
transform 1 0 88368 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_808
timestamp 1669390400
transform 1 0 91840 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_812
timestamp 1669390400
transform 1 0 92288 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_818
timestamp 1669390400
transform 1 0 92960 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_851
timestamp 1669390400
transform 1 0 96656 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_855
timestamp 1669390400
transform 1 0 97104 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_859
timestamp 1669390400
transform 1 0 97552 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_863
timestamp 1669390400
transform 1 0 98000 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_865
timestamp 1669390400
transform 1 0 98224 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_2
timestamp 1669390400
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_66
timestamp 1669390400
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_70
timestamp 1669390400
transform 1 0 9184 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1669390400
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_137
timestamp 1669390400
transform 1 0 16688 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1669390400
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_144
timestamp 1669390400
transform 1 0 17472 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_208
timestamp 1669390400
transform 1 0 24640 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1669390400
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1669390400
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_279
timestamp 1669390400
transform 1 0 32592 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1669390400
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1669390400
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_350
timestamp 1669390400
transform 1 0 40544 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1669390400
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1669390400
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_421
timestamp 1669390400
transform 1 0 48496 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1669390400
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_428
timestamp 1669390400
transform 1 0 49280 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_432
timestamp 1669390400
transform 1 0 49728 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_449
timestamp 1669390400
transform 1 0 51632 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_456
timestamp 1669390400
transform 1 0 52416 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_460
timestamp 1669390400
transform 1 0 52864 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_464
timestamp 1669390400
transform 1 0 53312 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_468
timestamp 1669390400
transform 1 0 53760 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_470
timestamp 1669390400
transform 1 0 53984 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_477
timestamp 1669390400
transform 1 0 54768 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_485
timestamp 1669390400
transform 1 0 55664 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_487
timestamp 1669390400
transform 1 0 55888 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_494
timestamp 1669390400
transform 1 0 56672 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1669390400
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_499
timestamp 1669390400
transform 1 0 57232 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_502
timestamp 1669390400
transform 1 0 57568 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_518
timestamp 1669390400
transform 1 0 59360 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_526
timestamp 1669390400
transform 1 0 60256 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_528
timestamp 1669390400
transform 1 0 60480 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_531
timestamp 1669390400
transform 1 0 60816 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_539
timestamp 1669390400
transform 1 0 61712 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_556
timestamp 1669390400
transform 1 0 63616 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_560
timestamp 1669390400
transform 1 0 64064 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_564
timestamp 1669390400
transform 1 0 64512 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_570
timestamp 1669390400
transform 1 0 65184 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_572
timestamp 1669390400
transform 1 0 65408 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_575
timestamp 1669390400
transform 1 0 65744 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_606
timestamp 1669390400
transform 1 0 69216 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_610
timestamp 1669390400
transform 1 0 69664 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_614
timestamp 1669390400
transform 1 0 70112 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_616
timestamp 1669390400
transform 1 0 70336 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_619
timestamp 1669390400
transform 1 0 70672 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_623
timestamp 1669390400
transform 1 0 71120 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_627
timestamp 1669390400
transform 1 0 71568 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_631
timestamp 1669390400
transform 1 0 72016 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_633
timestamp 1669390400
transform 1 0 72240 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_636
timestamp 1669390400
transform 1 0 72576 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1669390400
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_641
timestamp 1669390400
transform 1 0 73136 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_653
timestamp 1669390400
transform 1 0 74480 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_661
timestamp 1669390400
transform 1 0 75376 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_671
timestamp 1669390400
transform 1 0 76496 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_679
timestamp 1669390400
transform 1 0 77392 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_687
timestamp 1669390400
transform 1 0 78288 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_691
timestamp 1669390400
transform 1 0 78736 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_698
timestamp 1669390400
transform 1 0 79520 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_705
timestamp 1669390400
transform 1 0 80304 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_709
timestamp 1669390400
transform 1 0 80752 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_83_712
timestamp 1669390400
transform 1 0 81088 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_728
timestamp 1669390400
transform 1 0 82880 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_780
timestamp 1669390400
transform 1 0 88704 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_783
timestamp 1669390400
transform 1 0 89040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_799
timestamp 1669390400
transform 1 0 90832 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_851
timestamp 1669390400
transform 1 0 96656 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_854
timestamp 1669390400
transform 1 0 96992 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_83_862
timestamp 1669390400
transform 1 0 97888 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_2
timestamp 1669390400
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_34
timestamp 1669390400
transform 1 0 5152 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1669390400
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_101
timestamp 1669390400
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1669390400
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1669390400
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_172
timestamp 1669390400
transform 1 0 20608 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1669390400
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1669390400
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_243
timestamp 1669390400
transform 1 0 28560 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1669390400
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1669390400
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_314
timestamp 1669390400
transform 1 0 36512 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1669390400
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_321
timestamp 1669390400
transform 1 0 37296 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_385
timestamp 1669390400
transform 1 0 44464 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1669390400
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_392
timestamp 1669390400
transform 1 0 45248 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_424
timestamp 1669390400
transform 1 0 48832 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_428
timestamp 1669390400
transform 1 0 49280 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_458
timestamp 1669390400
transform 1 0 52640 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1669390400
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_463
timestamp 1669390400
transform 1 0 53200 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_494
timestamp 1669390400
transform 1 0 56672 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_525
timestamp 1669390400
transform 1 0 60144 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_529
timestamp 1669390400
transform 1 0 60592 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1669390400
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_534
timestamp 1669390400
transform 1 0 61152 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_585
timestamp 1669390400
transform 1 0 66864 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_589
timestamp 1669390400
transform 1 0 67312 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_595
timestamp 1669390400
transform 1 0 67984 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1669390400
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_605
timestamp 1669390400
transform 1 0 69104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_608
timestamp 1669390400
transform 1 0 69440 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_612
timestamp 1669390400
transform 1 0 69888 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_628
timestamp 1669390400
transform 1 0 71680 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_645
timestamp 1669390400
transform 1 0 73584 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_649
timestamp 1669390400
transform 1 0 74032 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_651
timestamp 1669390400
transform 1 0 74256 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_667
timestamp 1669390400
transform 1 0 76048 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_671
timestamp 1669390400
transform 1 0 76496 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1669390400
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_676
timestamp 1669390400
transform 1 0 77056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_692
timestamp 1669390400
transform 1 0 78848 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_696
timestamp 1669390400
transform 1 0 79296 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_700
timestamp 1669390400
transform 1 0 79744 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_704
timestamp 1669390400
transform 1 0 80192 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_712
timestamp 1669390400
transform 1 0 81088 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_715
timestamp 1669390400
transform 1 0 81424 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_723
timestamp 1669390400
transform 1 0 82320 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_725
timestamp 1669390400
transform 1 0 82544 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_728
timestamp 1669390400
transform 1 0 82880 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_735
timestamp 1669390400
transform 1 0 83664 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_744
timestamp 1669390400
transform 1 0 84672 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_747
timestamp 1669390400
transform 1 0 85008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_777
timestamp 1669390400
transform 1 0 88368 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_784
timestamp 1669390400
transform 1 0 89152 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_815
timestamp 1669390400
transform 1 0 92624 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_818
timestamp 1669390400
transform 1 0 92960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_825
timestamp 1669390400
transform 1 0 93744 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_829
timestamp 1669390400
transform 1 0 94192 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_833
timestamp 1669390400
transform 1 0 94640 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_863
timestamp 1669390400
transform 1 0 98000 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_865
timestamp 1669390400
transform 1 0 98224 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_2
timestamp 1669390400
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_66
timestamp 1669390400
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_70
timestamp 1669390400
transform 1 0 9184 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1669390400
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_137
timestamp 1669390400
transform 1 0 16688 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1669390400
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1669390400
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_208
timestamp 1669390400
transform 1 0 24640 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1669390400
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1669390400
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_279
timestamp 1669390400
transform 1 0 32592 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1669390400
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_286
timestamp 1669390400
transform 1 0 33376 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_350
timestamp 1669390400
transform 1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1669390400
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_357
timestamp 1669390400
transform 1 0 41328 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_421
timestamp 1669390400
transform 1 0 48496 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1669390400
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_428
timestamp 1669390400
transform 1 0 49280 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_444
timestamp 1669390400
transform 1 0 51072 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1669390400
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_499
timestamp 1669390400
transform 1 0 57232 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_515
timestamp 1669390400
transform 1 0 59024 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_519
timestamp 1669390400
transform 1 0 59472 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_523
timestamp 1669390400
transform 1 0 59920 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_556
timestamp 1669390400
transform 1 0 63616 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_560
timestamp 1669390400
transform 1 0 64064 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_570
timestamp 1669390400
transform 1 0 65184 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_574
timestamp 1669390400
transform 1 0 65632 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_576
timestamp 1669390400
transform 1 0 65856 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_592
timestamp 1669390400
transform 1 0 67648 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_594
timestamp 1669390400
transform 1 0 67872 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_624
timestamp 1669390400
transform 1 0 71232 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_628
timestamp 1669390400
transform 1 0 71680 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1669390400
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_641
timestamp 1669390400
transform 1 0 73136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_644
timestamp 1669390400
transform 1 0 73472 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_677
timestamp 1669390400
transform 1 0 77168 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_708
timestamp 1669390400
transform 1 0 80640 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_712
timestamp 1669390400
transform 1 0 81088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_715
timestamp 1669390400
transform 1 0 81424 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_752
timestamp 1669390400
transform 1 0 85568 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_760
timestamp 1669390400
transform 1 0 86464 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_764
timestamp 1669390400
transform 1 0 86912 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_768
timestamp 1669390400
transform 1 0 87360 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_772
timestamp 1669390400
transform 1 0 87808 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_776
timestamp 1669390400
transform 1 0 88256 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_780
timestamp 1669390400
transform 1 0 88704 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_783
timestamp 1669390400
transform 1 0 89040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_790
timestamp 1669390400
transform 1 0 89824 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_797
timestamp 1669390400
transform 1 0 90608 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_828
timestamp 1669390400
transform 1 0 94080 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_847
timestamp 1669390400
transform 1 0 96208 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_851
timestamp 1669390400
transform 1 0 96656 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_854
timestamp 1669390400
transform 1 0 96992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_857
timestamp 1669390400
transform 1 0 97328 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_865
timestamp 1669390400
transform 1 0 98224 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_2
timestamp 1669390400
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_34
timestamp 1669390400
transform 1 0 5152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1669390400
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_101
timestamp 1669390400
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1669390400
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1669390400
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_172
timestamp 1669390400
transform 1 0 20608 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1669390400
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1669390400
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_243
timestamp 1669390400
transform 1 0 28560 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1669390400
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_250
timestamp 1669390400
transform 1 0 29344 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_314
timestamp 1669390400
transform 1 0 36512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1669390400
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_321
timestamp 1669390400
transform 1 0 37296 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_385
timestamp 1669390400
transform 1 0 44464 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1669390400
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_392
timestamp 1669390400
transform 1 0 45248 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_408
timestamp 1669390400
transform 1 0 47040 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_412
timestamp 1669390400
transform 1 0 47488 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_420
timestamp 1669390400
transform 1 0 48384 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_451
timestamp 1669390400
transform 1 0 51856 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_455
timestamp 1669390400
transform 1 0 52304 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_457
timestamp 1669390400
transform 1 0 52528 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_460
timestamp 1669390400
transform 1 0 52864 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_463
timestamp 1669390400
transform 1 0 53200 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_471
timestamp 1669390400
transform 1 0 54096 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_475
timestamp 1669390400
transform 1 0 54544 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_477
timestamp 1669390400
transform 1 0 54768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_507
timestamp 1669390400
transform 1 0 58128 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_524
timestamp 1669390400
transform 1 0 60032 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_528
timestamp 1669390400
transform 1 0 60480 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_534
timestamp 1669390400
transform 1 0 61152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_564
timestamp 1669390400
transform 1 0 64512 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_568
timestamp 1669390400
transform 1 0 64960 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_576
timestamp 1669390400
transform 1 0 65856 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_578
timestamp 1669390400
transform 1 0 66080 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_585
timestamp 1669390400
transform 1 0 66864 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_587
timestamp 1669390400
transform 1 0 67088 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_590
timestamp 1669390400
transform 1 0 67424 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_594
timestamp 1669390400
transform 1 0 67872 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1669390400
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_605
timestamp 1669390400
transform 1 0 69104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_656
timestamp 1669390400
transform 1 0 74816 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_664
timestamp 1669390400
transform 1 0 75712 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_668
timestamp 1669390400
transform 1 0 76160 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_672
timestamp 1669390400
transform 1 0 76608 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_676
timestamp 1669390400
transform 1 0 77056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_679
timestamp 1669390400
transform 1 0 77392 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_683
timestamp 1669390400
transform 1 0 77840 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_699
timestamp 1669390400
transform 1 0 79632 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_703
timestamp 1669390400
transform 1 0 80080 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_707
timestamp 1669390400
transform 1 0 80528 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_711
timestamp 1669390400
transform 1 0 80976 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_713
timestamp 1669390400
transform 1 0 81200 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_716
timestamp 1669390400
transform 1 0 81536 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_733
timestamp 1669390400
transform 1 0 83440 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_737
timestamp 1669390400
transform 1 0 83888 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_741
timestamp 1669390400
transform 1 0 84336 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_744
timestamp 1669390400
transform 1 0 84672 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_747
timestamp 1669390400
transform 1 0 85008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_763
timestamp 1669390400
transform 1 0 86800 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_767
timestamp 1669390400
transform 1 0 87248 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_798
timestamp 1669390400
transform 1 0 90720 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_815
timestamp 1669390400
transform 1 0 92624 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_818
timestamp 1669390400
transform 1 0 92960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_821
timestamp 1669390400
transform 1 0 93296 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_825
timestamp 1669390400
transform 1 0 93744 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_829
timestamp 1669390400
transform 1 0 94192 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_839
timestamp 1669390400
transform 1 0 95312 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_847
timestamp 1669390400
transform 1 0 96208 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_851
timestamp 1669390400
transform 1 0 96656 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_859
timestamp 1669390400
transform 1 0 97552 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_863
timestamp 1669390400
transform 1 0 98000 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_865
timestamp 1669390400
transform 1 0 98224 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_2
timestamp 1669390400
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_66
timestamp 1669390400
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_70
timestamp 1669390400
transform 1 0 9184 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1669390400
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_137
timestamp 1669390400
transform 1 0 16688 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1669390400
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1669390400
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_208
timestamp 1669390400
transform 1 0 24640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1669390400
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1669390400
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_279
timestamp 1669390400
transform 1 0 32592 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1669390400
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_286
timestamp 1669390400
transform 1 0 33376 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_350
timestamp 1669390400
transform 1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1669390400
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_357
timestamp 1669390400
transform 1 0 41328 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_421
timestamp 1669390400
transform 1 0 48496 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1669390400
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_428
timestamp 1669390400
transform 1 0 49280 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_451
timestamp 1669390400
transform 1 0 51856 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_455
timestamp 1669390400
transform 1 0 52304 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_459
timestamp 1669390400
transform 1 0 52752 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_465
timestamp 1669390400
transform 1 0 53424 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_496
timestamp 1669390400
transform 1 0 56896 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_499
timestamp 1669390400
transform 1 0 57232 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_550
timestamp 1669390400
transform 1 0 62944 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_554
timestamp 1669390400
transform 1 0 63392 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_558
timestamp 1669390400
transform 1 0 63840 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_566
timestamp 1669390400
transform 1 0 64736 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_570
timestamp 1669390400
transform 1 0 65184 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_574
timestamp 1669390400
transform 1 0 65632 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_576
timestamp 1669390400
transform 1 0 65856 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_579
timestamp 1669390400
transform 1 0 66192 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_587
timestamp 1669390400
transform 1 0 67088 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_591
timestamp 1669390400
transform 1 0 67536 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_593
timestamp 1669390400
transform 1 0 67760 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_596
timestamp 1669390400
transform 1 0 68096 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_598
timestamp 1669390400
transform 1 0 68320 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_605
timestamp 1669390400
transform 1 0 69104 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_636
timestamp 1669390400
transform 1 0 72576 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_638
timestamp 1669390400
transform 1 0 72800 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_641
timestamp 1669390400
transform 1 0 73136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_644
timestamp 1669390400
transform 1 0 73472 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_654
timestamp 1669390400
transform 1 0 74592 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_658
timestamp 1669390400
transform 1 0 75040 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_662
timestamp 1669390400
transform 1 0 75488 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_666
timestamp 1669390400
transform 1 0 75936 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_670
timestamp 1669390400
transform 1 0 76384 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_674
timestamp 1669390400
transform 1 0 76832 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_678
timestamp 1669390400
transform 1 0 77280 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_709
timestamp 1669390400
transform 1 0 80752 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_712
timestamp 1669390400
transform 1 0 81088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_742
timestamp 1669390400
transform 1 0 84448 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_774
timestamp 1669390400
transform 1 0 88032 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_778
timestamp 1669390400
transform 1 0 88480 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_780
timestamp 1669390400
transform 1 0 88704 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_783
timestamp 1669390400
transform 1 0 89040 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_787
timestamp 1669390400
transform 1 0 89488 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_839
timestamp 1669390400
transform 1 0 95312 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_843
timestamp 1669390400
transform 1 0 95760 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_851
timestamp 1669390400
transform 1 0 96656 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_87_854
timestamp 1669390400
transform 1 0 96992 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_862
timestamp 1669390400
transform 1 0 97888 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_2
timestamp 1669390400
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1669390400
transform 1 0 5152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1669390400
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_101
timestamp 1669390400
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1669390400
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1669390400
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_172
timestamp 1669390400
transform 1 0 20608 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1669390400
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1669390400
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_243
timestamp 1669390400
transform 1 0 28560 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1669390400
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_250
timestamp 1669390400
transform 1 0 29344 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_314
timestamp 1669390400
transform 1 0 36512 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1669390400
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_321
timestamp 1669390400
transform 1 0 37296 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_385
timestamp 1669390400
transform 1 0 44464 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_389
timestamp 1669390400
transform 1 0 44912 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_392
timestamp 1669390400
transform 1 0 45248 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_424
timestamp 1669390400
transform 1 0 48832 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_428
timestamp 1669390400
transform 1 0 49280 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_436
timestamp 1669390400
transform 1 0 50176 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_452
timestamp 1669390400
transform 1 0 51968 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1669390400
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_463
timestamp 1669390400
transform 1 0 53200 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_471
timestamp 1669390400
transform 1 0 54096 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_477
timestamp 1669390400
transform 1 0 54768 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_485
timestamp 1669390400
transform 1 0 55664 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_502
timestamp 1669390400
transform 1 0 57568 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_519
timestamp 1669390400
transform 1 0 59472 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_523
timestamp 1669390400
transform 1 0 59920 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_531
timestamp 1669390400
transform 1 0 60816 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_534
timestamp 1669390400
transform 1 0 61152 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_536
timestamp 1669390400
transform 1 0 61376 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_552
timestamp 1669390400
transform 1 0 63168 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_569
timestamp 1669390400
transform 1 0 65072 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_573
timestamp 1669390400
transform 1 0 65520 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_577
timestamp 1669390400
transform 1 0 65968 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_593
timestamp 1669390400
transform 1 0 67760 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_601
timestamp 1669390400
transform 1 0 68656 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_605
timestamp 1669390400
transform 1 0 69104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_608
timestamp 1669390400
transform 1 0 69440 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_622
timestamp 1669390400
transform 1 0 71008 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_626
timestamp 1669390400
transform 1 0 71456 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_635
timestamp 1669390400
transform 1 0 72464 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_639
timestamp 1669390400
transform 1 0 72912 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_641
timestamp 1669390400
transform 1 0 73136 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_650
timestamp 1669390400
transform 1 0 74144 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_669
timestamp 1669390400
transform 1 0 76272 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_673
timestamp 1669390400
transform 1 0 76720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_676
timestamp 1669390400
transform 1 0 77056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_679
timestamp 1669390400
transform 1 0 77392 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_681
timestamp 1669390400
transform 1 0 77616 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_684
timestamp 1669390400
transform 1 0 77952 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_688
timestamp 1669390400
transform 1 0 78400 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_740
timestamp 1669390400
transform 1 0 84224 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_744
timestamp 1669390400
transform 1 0 84672 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_747
timestamp 1669390400
transform 1 0 85008 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_755
timestamp 1669390400
transform 1 0 85904 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_759
timestamp 1669390400
transform 1 0 86352 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_763
timestamp 1669390400
transform 1 0 86800 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_815
timestamp 1669390400
transform 1 0 92624 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_818
timestamp 1669390400
transform 1 0 92960 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_826
timestamp 1669390400
transform 1 0 93856 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_830
timestamp 1669390400
transform 1 0 94304 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_863
timestamp 1669390400
transform 1 0 98000 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_865
timestamp 1669390400
transform 1 0 98224 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_2
timestamp 1669390400
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_66
timestamp 1669390400
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_70
timestamp 1669390400
transform 1 0 9184 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1669390400
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_137
timestamp 1669390400
transform 1 0 16688 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1669390400
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1669390400
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_208
timestamp 1669390400
transform 1 0 24640 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1669390400
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_215
timestamp 1669390400
transform 1 0 25424 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_279
timestamp 1669390400
transform 1 0 32592 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1669390400
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_286
timestamp 1669390400
transform 1 0 33376 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_350
timestamp 1669390400
transform 1 0 40544 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1669390400
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_357
timestamp 1669390400
transform 1 0 41328 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_421
timestamp 1669390400
transform 1 0 48496 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1669390400
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_428
timestamp 1669390400
transform 1 0 49280 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_444
timestamp 1669390400
transform 1 0 51072 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_448
timestamp 1669390400
transform 1 0 51520 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_450
timestamp 1669390400
transform 1 0 51744 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_453
timestamp 1669390400
transform 1 0 52080 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_485
timestamp 1669390400
transform 1 0 55664 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_493
timestamp 1669390400
transform 1 0 56560 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_499
timestamp 1669390400
transform 1 0 57232 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_502
timestamp 1669390400
transform 1 0 57568 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_506
timestamp 1669390400
transform 1 0 58016 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_510
timestamp 1669390400
transform 1 0 58464 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_518
timestamp 1669390400
transform 1 0 59360 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_521
timestamp 1669390400
transform 1 0 59696 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_529
timestamp 1669390400
transform 1 0 60592 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_533
timestamp 1669390400
transform 1 0 61040 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_564
timestamp 1669390400
transform 1 0 64512 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_570
timestamp 1669390400
transform 1 0 65184 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_573
timestamp 1669390400
transform 1 0 65520 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_589
timestamp 1669390400
transform 1 0 67312 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_593
timestamp 1669390400
transform 1 0 67760 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_595
timestamp 1669390400
transform 1 0 67984 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_602
timestamp 1669390400
transform 1 0 68768 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_618
timestamp 1669390400
transform 1 0 70560 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_622
timestamp 1669390400
transform 1 0 71008 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_625
timestamp 1669390400
transform 1 0 71344 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_633
timestamp 1669390400
transform 1 0 72240 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_637
timestamp 1669390400
transform 1 0 72688 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_641
timestamp 1669390400
transform 1 0 73136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_644
timestamp 1669390400
transform 1 0 73472 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_648
timestamp 1669390400
transform 1 0 73920 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_679
timestamp 1669390400
transform 1 0 77392 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_683
timestamp 1669390400
transform 1 0 77840 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_699
timestamp 1669390400
transform 1 0 79632 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_703
timestamp 1669390400
transform 1 0 80080 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_707
timestamp 1669390400
transform 1 0 80528 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_709
timestamp 1669390400
transform 1 0 80752 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_712
timestamp 1669390400
transform 1 0 81088 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_720
timestamp 1669390400
transform 1 0 81984 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_724
timestamp 1669390400
transform 1 0 82432 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_726
timestamp 1669390400
transform 1 0 82656 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_89_733
timestamp 1669390400
transform 1 0 83440 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_765
timestamp 1669390400
transform 1 0 87024 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_773
timestamp 1669390400
transform 1 0 87920 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_780
timestamp 1669390400
transform 1 0 88704 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_783
timestamp 1669390400
transform 1 0 89040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_799
timestamp 1669390400
transform 1 0 90832 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_803
timestamp 1669390400
transform 1 0 91280 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_89_811
timestamp 1669390400
transform 1 0 92176 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_819
timestamp 1669390400
transform 1 0 93072 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_823
timestamp 1669390400
transform 1 0 93520 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_826
timestamp 1669390400
transform 1 0 93856 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_830
timestamp 1669390400
transform 1 0 94304 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_834
timestamp 1669390400
transform 1 0 94752 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_851
timestamp 1669390400
transform 1 0 96656 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_854
timestamp 1669390400
transform 1 0 96992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_861
timestamp 1669390400
transform 1 0 97776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_865
timestamp 1669390400
transform 1 0 98224 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_2
timestamp 1669390400
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_34
timestamp 1669390400
transform 1 0 5152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1669390400
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_101
timestamp 1669390400
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1669390400
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1669390400
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_172
timestamp 1669390400
transform 1 0 20608 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1669390400
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1669390400
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_243
timestamp 1669390400
transform 1 0 28560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1669390400
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_250
timestamp 1669390400
transform 1 0 29344 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_314
timestamp 1669390400
transform 1 0 36512 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1669390400
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_321
timestamp 1669390400
transform 1 0 37296 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_385
timestamp 1669390400
transform 1 0 44464 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1669390400
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_392
timestamp 1669390400
transform 1 0 45248 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_424
timestamp 1669390400
transform 1 0 48832 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_432
timestamp 1669390400
transform 1 0 49728 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_434
timestamp 1669390400
transform 1 0 49952 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_437
timestamp 1669390400
transform 1 0 50288 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_444
timestamp 1669390400
transform 1 0 51072 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_451
timestamp 1669390400
transform 1 0 51856 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_458
timestamp 1669390400
transform 1 0 52640 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_460
timestamp 1669390400
transform 1 0 52864 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_463
timestamp 1669390400
transform 1 0 53200 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_466
timestamp 1669390400
transform 1 0 53536 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_470
timestamp 1669390400
transform 1 0 53984 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_474
timestamp 1669390400
transform 1 0 54432 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_478
timestamp 1669390400
transform 1 0 54880 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_510
timestamp 1669390400
transform 1 0 58464 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_518
timestamp 1669390400
transform 1 0 59360 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_520
timestamp 1669390400
transform 1 0 59584 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_523
timestamp 1669390400
transform 1 0 59920 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1669390400
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_534
timestamp 1669390400
transform 1 0 61152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_550
timestamp 1669390400
transform 1 0 62944 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_602
timestamp 1669390400
transform 1 0 68768 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_605
timestamp 1669390400
transform 1 0 69104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_621
timestamp 1669390400
transform 1 0 70896 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_625
timestamp 1669390400
transform 1 0 71344 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_635
timestamp 1669390400
transform 1 0 72464 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_639
timestamp 1669390400
transform 1 0 72912 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_647
timestamp 1669390400
transform 1 0 73808 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_651
timestamp 1669390400
transform 1 0 74256 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_653
timestamp 1669390400
transform 1 0 74480 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_660
timestamp 1669390400
transform 1 0 75264 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_664
timestamp 1669390400
transform 1 0 75712 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_673
timestamp 1669390400
transform 1 0 76720 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_676
timestamp 1669390400
transform 1 0 77056 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_678
timestamp 1669390400
transform 1 0 77280 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_681
timestamp 1669390400
transform 1 0 77616 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_691
timestamp 1669390400
transform 1 0 78736 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_707
timestamp 1669390400
transform 1 0 80528 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_715
timestamp 1669390400
transform 1 0 81424 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_719
timestamp 1669390400
transform 1 0 81872 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_723
timestamp 1669390400
transform 1 0 82320 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_727
timestamp 1669390400
transform 1 0 82768 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_734
timestamp 1669390400
transform 1 0 83552 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_738
timestamp 1669390400
transform 1 0 84000 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_742
timestamp 1669390400
transform 1 0 84448 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_744
timestamp 1669390400
transform 1 0 84672 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_747
timestamp 1669390400
transform 1 0 85008 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_90_763
timestamp 1669390400
transform 1 0 86800 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_800
timestamp 1669390400
transform 1 0 90944 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_804
timestamp 1669390400
transform 1 0 91392 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_808
timestamp 1669390400
transform 1 0 91840 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_812
timestamp 1669390400
transform 1 0 92288 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_818
timestamp 1669390400
transform 1 0 92960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_821
timestamp 1669390400
transform 1 0 93296 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_825
timestamp 1669390400
transform 1 0 93744 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_829
timestamp 1669390400
transform 1 0 94192 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_833
timestamp 1669390400
transform 1 0 94640 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_863
timestamp 1669390400
transform 1 0 98000 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_865
timestamp 1669390400
transform 1 0 98224 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_2
timestamp 1669390400
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_66
timestamp 1669390400
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_70
timestamp 1669390400
transform 1 0 9184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1669390400
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_137
timestamp 1669390400
transform 1 0 16688 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1669390400
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1669390400
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_208
timestamp 1669390400
transform 1 0 24640 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1669390400
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_215
timestamp 1669390400
transform 1 0 25424 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_279
timestamp 1669390400
transform 1 0 32592 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1669390400
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_286
timestamp 1669390400
transform 1 0 33376 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_350
timestamp 1669390400
transform 1 0 40544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1669390400
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_357
timestamp 1669390400
transform 1 0 41328 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_421
timestamp 1669390400
transform 1 0 48496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1669390400
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_428
timestamp 1669390400
transform 1 0 49280 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_432
timestamp 1669390400
transform 1 0 49728 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_462
timestamp 1669390400
transform 1 0 53088 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_469
timestamp 1669390400
transform 1 0 53872 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_476
timestamp 1669390400
transform 1 0 54656 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_483
timestamp 1669390400
transform 1 0 55440 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_490
timestamp 1669390400
transform 1 0 56224 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_494
timestamp 1669390400
transform 1 0 56672 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1669390400
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_499
timestamp 1669390400
transform 1 0 57232 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_502
timestamp 1669390400
transform 1 0 57568 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_506
timestamp 1669390400
transform 1 0 58016 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_522
timestamp 1669390400
transform 1 0 59808 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_526
timestamp 1669390400
transform 1 0 60256 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_556
timestamp 1669390400
transform 1 0 63616 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_560
timestamp 1669390400
transform 1 0 64064 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_564
timestamp 1669390400
transform 1 0 64512 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_570
timestamp 1669390400
transform 1 0 65184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_577
timestamp 1669390400
transform 1 0 65968 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_581
timestamp 1669390400
transform 1 0 66416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_614
timestamp 1669390400
transform 1 0 70112 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_631
timestamp 1669390400
transform 1 0 72016 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_635
timestamp 1669390400
transform 1 0 72464 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_641
timestamp 1669390400
transform 1 0 73136 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_645
timestamp 1669390400
transform 1 0 73584 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_648
timestamp 1669390400
transform 1 0 73920 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_656
timestamp 1669390400
transform 1 0 74816 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_660
timestamp 1669390400
transform 1 0 75264 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_662
timestamp 1669390400
transform 1 0 75488 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_665
timestamp 1669390400
transform 1 0 75824 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_669
timestamp 1669390400
transform 1 0 76272 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_701
timestamp 1669390400
transform 1 0 79856 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_709
timestamp 1669390400
transform 1 0 80752 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_712
timestamp 1669390400
transform 1 0 81088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_715
timestamp 1669390400
transform 1 0 81424 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_746
timestamp 1669390400
transform 1 0 84896 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_750
timestamp 1669390400
transform 1 0 85344 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_766
timestamp 1669390400
transform 1 0 87136 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_780
timestamp 1669390400
transform 1 0 88704 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_783
timestamp 1669390400
transform 1 0 89040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_799
timestamp 1669390400
transform 1 0 90832 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_801
timestamp 1669390400
transform 1 0 91056 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_817
timestamp 1669390400
transform 1 0 92848 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_819
timestamp 1669390400
transform 1 0 93072 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_835
timestamp 1669390400
transform 1 0 94864 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_839
timestamp 1669390400
transform 1 0 95312 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_846
timestamp 1669390400
transform 1 0 96096 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_850
timestamp 1669390400
transform 1 0 96544 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_854
timestamp 1669390400
transform 1 0 96992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_857
timestamp 1669390400
transform 1 0 97328 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_865
timestamp 1669390400
transform 1 0 98224 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_2
timestamp 1669390400
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_34
timestamp 1669390400
transform 1 0 5152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1669390400
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1669390400
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1669390400
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_108
timestamp 1669390400
transform 1 0 13440 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_172
timestamp 1669390400
transform 1 0 20608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1669390400
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_179
timestamp 1669390400
transform 1 0 21392 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_243
timestamp 1669390400
transform 1 0 28560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1669390400
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_250
timestamp 1669390400
transform 1 0 29344 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_314
timestamp 1669390400
transform 1 0 36512 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1669390400
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_321
timestamp 1669390400
transform 1 0 37296 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_385
timestamp 1669390400
transform 1 0 44464 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_389
timestamp 1669390400
transform 1 0 44912 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_92_392
timestamp 1669390400
transform 1 0 45248 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_424
timestamp 1669390400
transform 1 0 48832 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_428
timestamp 1669390400
transform 1 0 49280 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_430
timestamp 1669390400
transform 1 0 49504 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_460
timestamp 1669390400
transform 1 0 52864 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_463
timestamp 1669390400
transform 1 0 53200 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_496
timestamp 1669390400
transform 1 0 56896 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_527
timestamp 1669390400
transform 1 0 60368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1669390400
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_534
timestamp 1669390400
transform 1 0 61152 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_548
timestamp 1669390400
transform 1 0 62720 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_552
timestamp 1669390400
transform 1 0 63168 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_585
timestamp 1669390400
transform 1 0 66864 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_589
timestamp 1669390400
transform 1 0 67312 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_593
timestamp 1669390400
transform 1 0 67760 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_597
timestamp 1669390400
transform 1 0 68208 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_601
timestamp 1669390400
transform 1 0 68656 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_605
timestamp 1669390400
transform 1 0 69104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_612
timestamp 1669390400
transform 1 0 69888 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_616
timestamp 1669390400
transform 1 0 70336 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_620
timestamp 1669390400
transform 1 0 70784 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_626
timestamp 1669390400
transform 1 0 71456 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_644
timestamp 1669390400
transform 1 0 73472 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_648
timestamp 1669390400
transform 1 0 73920 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_655
timestamp 1669390400
transform 1 0 74704 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_663
timestamp 1669390400
transform 1 0 75600 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_670
timestamp 1669390400
transform 1 0 76384 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_676
timestamp 1669390400
transform 1 0 77056 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_721
timestamp 1669390400
transform 1 0 82096 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_728
timestamp 1669390400
transform 1 0 82880 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_735
timestamp 1669390400
transform 1 0 83664 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_744
timestamp 1669390400
transform 1 0 84672 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_747
timestamp 1669390400
transform 1 0 85008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_753
timestamp 1669390400
transform 1 0 85680 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_760
timestamp 1669390400
transform 1 0 86464 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_92_764
timestamp 1669390400
transform 1 0 86912 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_780
timestamp 1669390400
transform 1 0 88704 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_784
timestamp 1669390400
transform 1 0 89152 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_815
timestamp 1669390400
transform 1 0 92624 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_818
timestamp 1669390400
transform 1 0 92960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_848
timestamp 1669390400
transform 1 0 96320 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_865
timestamp 1669390400
transform 1 0 98224 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_2
timestamp 1669390400
transform 1 0 1568 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_66
timestamp 1669390400
transform 1 0 8736 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_70
timestamp 1669390400
transform 1 0 9184 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_73
timestamp 1669390400
transform 1 0 9520 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_137
timestamp 1669390400
transform 1 0 16688 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_141
timestamp 1669390400
transform 1 0 17136 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_144
timestamp 1669390400
transform 1 0 17472 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_208
timestamp 1669390400
transform 1 0 24640 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_212
timestamp 1669390400
transform 1 0 25088 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_215
timestamp 1669390400
transform 1 0 25424 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_279
timestamp 1669390400
transform 1 0 32592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_283
timestamp 1669390400
transform 1 0 33040 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_286
timestamp 1669390400
transform 1 0 33376 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_350
timestamp 1669390400
transform 1 0 40544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_354
timestamp 1669390400
transform 1 0 40992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_93_357
timestamp 1669390400
transform 1 0 41328 0 -1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_421
timestamp 1669390400
transform 1 0 48496 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_425
timestamp 1669390400
transform 1 0 48944 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_428
timestamp 1669390400
transform 1 0 49280 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_436
timestamp 1669390400
transform 1 0 50176 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_440
timestamp 1669390400
transform 1 0 50624 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_444
timestamp 1669390400
transform 1 0 51072 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_496
timestamp 1669390400
transform 1 0 56896 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_499
timestamp 1669390400
transform 1 0 57232 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_505
timestamp 1669390400
transform 1 0 57904 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_512
timestamp 1669390400
transform 1 0 58688 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_93_516
timestamp 1669390400
transform 1 0 59136 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_548
timestamp 1669390400
transform 1 0 62720 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_552
timestamp 1669390400
transform 1 0 63168 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_556
timestamp 1669390400
transform 1 0 63616 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_560
timestamp 1669390400
transform 1 0 64064 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_567
timestamp 1669390400
transform 1 0 64848 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_570
timestamp 1669390400
transform 1 0 65184 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_577
timestamp 1669390400
transform 1 0 65968 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_584
timestamp 1669390400
transform 1 0 66752 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_591
timestamp 1669390400
transform 1 0 67536 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_624
timestamp 1669390400
transform 1 0 71232 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_634
timestamp 1669390400
transform 1 0 72352 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_638
timestamp 1669390400
transform 1 0 72800 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_641
timestamp 1669390400
transform 1 0 73136 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_643
timestamp 1669390400
transform 1 0 73360 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_673
timestamp 1669390400
transform 1 0 76720 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_677
timestamp 1669390400
transform 1 0 77168 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_681
timestamp 1669390400
transform 1 0 77616 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_684
timestamp 1669390400
transform 1 0 77952 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_688
timestamp 1669390400
transform 1 0 78400 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_691
timestamp 1669390400
transform 1 0 78736 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_699
timestamp 1669390400
transform 1 0 79632 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_705
timestamp 1669390400
transform 1 0 80304 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_709
timestamp 1669390400
transform 1 0 80752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_712
timestamp 1669390400
transform 1 0 81088 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_718
timestamp 1669390400
transform 1 0 81760 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_725
timestamp 1669390400
transform 1 0 82544 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_729
timestamp 1669390400
transform 1 0 82992 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_731
timestamp 1669390400
transform 1 0 83216 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_761
timestamp 1669390400
transform 1 0 86576 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_768
timestamp 1669390400
transform 1 0 87360 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_772
timestamp 1669390400
transform 1 0 87808 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_780
timestamp 1669390400
transform 1 0 88704 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_783
timestamp 1669390400
transform 1 0 89040 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_791
timestamp 1669390400
transform 1 0 89936 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_799
timestamp 1669390400
transform 1 0 90832 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_851
timestamp 1669390400
transform 1 0 96656 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_854
timestamp 1669390400
transform 1 0 96992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_857
timestamp 1669390400
transform 1 0 97328 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_865
timestamp 1669390400
transform 1 0 98224 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_94_2
timestamp 1669390400
transform 1 0 1568 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_34
timestamp 1669390400
transform 1 0 5152 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_37
timestamp 1669390400
transform 1 0 5488 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_101
timestamp 1669390400
transform 1 0 12656 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_105
timestamp 1669390400
transform 1 0 13104 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_108
timestamp 1669390400
transform 1 0 13440 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_172
timestamp 1669390400
transform 1 0 20608 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_176
timestamp 1669390400
transform 1 0 21056 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_179
timestamp 1669390400
transform 1 0 21392 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_243
timestamp 1669390400
transform 1 0 28560 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_247
timestamp 1669390400
transform 1 0 29008 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_250
timestamp 1669390400
transform 1 0 29344 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_314
timestamp 1669390400
transform 1 0 36512 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_318
timestamp 1669390400
transform 1 0 36960 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_94_321
timestamp 1669390400
transform 1 0 37296 0 1 76832
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_385
timestamp 1669390400
transform 1 0 44464 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_389
timestamp 1669390400
transform 1 0 44912 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_94_392
timestamp 1669390400
transform 1 0 45248 0 1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_424
timestamp 1669390400
transform 1 0 48832 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_428
timestamp 1669390400
transform 1 0 49280 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_430
timestamp 1669390400
transform 1 0 49504 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_460
timestamp 1669390400
transform 1 0 52864 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_463
timestamp 1669390400
transform 1 0 53200 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_466
timestamp 1669390400
transform 1 0 53536 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_470
timestamp 1669390400
transform 1 0 53984 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_501
timestamp 1669390400
transform 1 0 57456 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_505
timestamp 1669390400
transform 1 0 57904 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_509
timestamp 1669390400
transform 1 0 58352 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_513
timestamp 1669390400
transform 1 0 58800 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_529
timestamp 1669390400
transform 1 0 60592 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_531
timestamp 1669390400
transform 1 0 60816 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_534
timestamp 1669390400
transform 1 0 61152 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_544
timestamp 1669390400
transform 1 0 62272 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_596
timestamp 1669390400
transform 1 0 68096 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_600
timestamp 1669390400
transform 1 0 68544 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_602
timestamp 1669390400
transform 1 0 68768 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_605
timestamp 1669390400
transform 1 0 69104 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_608
timestamp 1669390400
transform 1 0 69440 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_612
timestamp 1669390400
transform 1 0 69888 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_622
timestamp 1669390400
transform 1 0 71008 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_626
timestamp 1669390400
transform 1 0 71456 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_633
timestamp 1669390400
transform 1 0 72240 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_635
timestamp 1669390400
transform 1 0 72464 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_641
timestamp 1669390400
transform 1 0 73136 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_649
timestamp 1669390400
transform 1 0 74032 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_652
timestamp 1669390400
transform 1 0 74368 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_659
timestamp 1669390400
transform 1 0 75152 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_667
timestamp 1669390400
transform 1 0 76048 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_673
timestamp 1669390400
transform 1 0 76720 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_676
timestamp 1669390400
transform 1 0 77056 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_682
timestamp 1669390400
transform 1 0 77728 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_689
timestamp 1669390400
transform 1 0 78512 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_697
timestamp 1669390400
transform 1 0 79408 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_703
timestamp 1669390400
transform 1 0 80080 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_707
timestamp 1669390400
transform 1 0 80528 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_711
timestamp 1669390400
transform 1 0 80976 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_720
timestamp 1669390400
transform 1 0 81984 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_724
timestamp 1669390400
transform 1 0 82432 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_733
timestamp 1669390400
transform 1 0 83440 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_737
timestamp 1669390400
transform 1 0 83888 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_743
timestamp 1669390400
transform 1 0 84560 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_747
timestamp 1669390400
transform 1 0 85008 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_777
timestamp 1669390400
transform 1 0 88368 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_781
timestamp 1669390400
transform 1 0 88816 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_797
timestamp 1669390400
transform 1 0 90608 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_801
timestamp 1669390400
transform 1 0 91056 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_809
timestamp 1669390400
transform 1 0 91952 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_815
timestamp 1669390400
transform 1 0 92624 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_818
timestamp 1669390400
transform 1 0 92960 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_825
timestamp 1669390400
transform 1 0 93744 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_829
timestamp 1669390400
transform 1 0 94192 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_94_831
timestamp 1669390400
transform 1 0 94416 0 1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_94_834
timestamp 1669390400
transform 1 0 94752 0 1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_94_838
timestamp 1669390400
transform 1 0 95200 0 1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_94_854
timestamp 1669390400
transform 1 0 96992 0 1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_94_862
timestamp 1669390400
transform 1 0 97888 0 1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_2
timestamp 1669390400
transform 1 0 1568 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_66
timestamp 1669390400
transform 1 0 8736 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_70
timestamp 1669390400
transform 1 0 9184 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_73
timestamp 1669390400
transform 1 0 9520 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_137
timestamp 1669390400
transform 1 0 16688 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_141
timestamp 1669390400
transform 1 0 17136 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_144
timestamp 1669390400
transform 1 0 17472 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_208
timestamp 1669390400
transform 1 0 24640 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_212
timestamp 1669390400
transform 1 0 25088 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_215
timestamp 1669390400
transform 1 0 25424 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_279
timestamp 1669390400
transform 1 0 32592 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_283
timestamp 1669390400
transform 1 0 33040 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_95_286
timestamp 1669390400
transform 1 0 33376 0 -1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_350
timestamp 1669390400
transform 1 0 40544 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_354
timestamp 1669390400
transform 1 0 40992 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_95_357
timestamp 1669390400
transform 1 0 41328 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_95_389
timestamp 1669390400
transform 1 0 44912 0 -1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_405
timestamp 1669390400
transform 1 0 46704 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_413
timestamp 1669390400
transform 1 0 47600 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_417
timestamp 1669390400
transform 1 0 48048 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_421
timestamp 1669390400
transform 1 0 48496 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_425
timestamp 1669390400
transform 1 0 48944 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_428
timestamp 1669390400
transform 1 0 49280 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_435
timestamp 1669390400
transform 1 0 50064 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_442
timestamp 1669390400
transform 1 0 50848 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_449
timestamp 1669390400
transform 1 0 51632 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_456
timestamp 1669390400
transform 1 0 52416 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_460
timestamp 1669390400
transform 1 0 52864 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_464
timestamp 1669390400
transform 1 0 53312 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_468
timestamp 1669390400
transform 1 0 53760 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_472
timestamp 1669390400
transform 1 0 54208 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_481
timestamp 1669390400
transform 1 0 55216 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_489
timestamp 1669390400
transform 1 0 56112 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_496
timestamp 1669390400
transform 1 0 56896 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_499
timestamp 1669390400
transform 1 0 57232 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_502
timestamp 1669390400
transform 1 0 57568 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_509
timestamp 1669390400
transform 1 0 58352 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_513
timestamp 1669390400
transform 1 0 58800 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_515
timestamp 1669390400
transform 1 0 59024 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_548
timestamp 1669390400
transform 1 0 62720 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_552
timestamp 1669390400
transform 1 0 63168 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_556
timestamp 1669390400
transform 1 0 63616 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_564
timestamp 1669390400
transform 1 0 64512 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_570
timestamp 1669390400
transform 1 0 65184 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_576
timestamp 1669390400
transform 1 0 65856 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_583
timestamp 1669390400
transform 1 0 66640 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_587
timestamp 1669390400
transform 1 0 67088 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_597
timestamp 1669390400
transform 1 0 68208 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_601
timestamp 1669390400
transform 1 0 68656 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_609
timestamp 1669390400
transform 1 0 69552 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_616
timestamp 1669390400
transform 1 0 70336 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_620
timestamp 1669390400
transform 1 0 70784 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_624
timestamp 1669390400
transform 1 0 71232 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_634
timestamp 1669390400
transform 1 0 72352 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_638
timestamp 1669390400
transform 1 0 72800 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_641
timestamp 1669390400
transform 1 0 73136 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_644
timestamp 1669390400
transform 1 0 73472 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_675
timestamp 1669390400
transform 1 0 76944 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_709
timestamp 1669390400
transform 1 0 80752 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_712
timestamp 1669390400
transform 1 0 81088 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_742
timestamp 1669390400
transform 1 0 84448 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_746
timestamp 1669390400
transform 1 0 84896 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_779
timestamp 1669390400
transform 1 0 88592 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_783
timestamp 1669390400
transform 1 0 89040 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_789
timestamp 1669390400
transform 1 0 89712 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_797
timestamp 1669390400
transform 1 0 90608 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_95_801
timestamp 1669390400
transform 1 0 91056 0 -1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_832
timestamp 1669390400
transform 1 0 94528 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_95_851
timestamp 1669390400
transform 1 0 96656 0 -1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_95_854
timestamp 1669390400
transform 1 0 96992 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_95_862
timestamp 1669390400
transform 1 0 97888 0 -1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_96_2
timestamp 1669390400
transform 1 0 1568 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_34
timestamp 1669390400
transform 1 0 5152 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_37
timestamp 1669390400
transform 1 0 5488 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_101
timestamp 1669390400
transform 1 0 12656 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_105
timestamp 1669390400
transform 1 0 13104 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_108
timestamp 1669390400
transform 1 0 13440 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_172
timestamp 1669390400
transform 1 0 20608 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_176
timestamp 1669390400
transform 1 0 21056 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_179
timestamp 1669390400
transform 1 0 21392 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_243
timestamp 1669390400
transform 1 0 28560 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_247
timestamp 1669390400
transform 1 0 29008 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_250
timestamp 1669390400
transform 1 0 29344 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_314
timestamp 1669390400
transform 1 0 36512 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_318
timestamp 1669390400
transform 1 0 36960 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_96_321
timestamp 1669390400
transform 1 0 37296 0 1 78400
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_385
timestamp 1669390400
transform 1 0 44464 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_389
timestamp 1669390400
transform 1 0 44912 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_96_392
timestamp 1669390400
transform 1 0 45248 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_424
timestamp 1669390400
transform 1 0 48832 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_426
timestamp 1669390400
transform 1 0 49056 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_429
timestamp 1669390400
transform 1 0 49392 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_433
timestamp 1669390400
transform 1 0 49840 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_437
timestamp 1669390400
transform 1 0 50288 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_444
timestamp 1669390400
transform 1 0 51072 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_451
timestamp 1669390400
transform 1 0 51856 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_458
timestamp 1669390400
transform 1 0 52640 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_460
timestamp 1669390400
transform 1 0 52864 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_463
timestamp 1669390400
transform 1 0 53200 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_469
timestamp 1669390400
transform 1 0 53872 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_473
timestamp 1669390400
transform 1 0 54320 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_96_477
timestamp 1669390400
transform 1 0 54768 0 1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_493
timestamp 1669390400
transform 1 0 56560 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_497
timestamp 1669390400
transform 1 0 57008 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_531
timestamp 1669390400
transform 1 0 60816 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_534
timestamp 1669390400
transform 1 0 61152 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_537
timestamp 1669390400
transform 1 0 61488 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_541
timestamp 1669390400
transform 1 0 61936 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_545
timestamp 1669390400
transform 1 0 62384 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_96_549
timestamp 1669390400
transform 1 0 62832 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_557
timestamp 1669390400
transform 1 0 63728 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_590
timestamp 1669390400
transform 1 0 67424 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_597
timestamp 1669390400
transform 1 0 68208 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_601
timestamp 1669390400
transform 1 0 68656 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_605
timestamp 1669390400
transform 1 0 69104 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_656
timestamp 1669390400
transform 1 0 74816 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_664
timestamp 1669390400
transform 1 0 75712 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_671
timestamp 1669390400
transform 1 0 76496 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_673
timestamp 1669390400
transform 1 0 76720 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_676
timestamp 1669390400
transform 1 0 77056 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_727
timestamp 1669390400
transform 1 0 82768 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_734
timestamp 1669390400
transform 1 0 83552 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_741
timestamp 1669390400
transform 1 0 84336 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_747
timestamp 1669390400
transform 1 0 85008 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_780
timestamp 1669390400
transform 1 0 88704 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_784
timestamp 1669390400
transform 1 0 89152 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_96_788
timestamp 1669390400
transform 1 0 89600 0 1 78400
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_96_810
timestamp 1669390400
transform 1 0 92064 0 1 78400
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_814
timestamp 1669390400
transform 1 0 92512 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_818
timestamp 1669390400
transform 1 0 92960 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_96_825
timestamp 1669390400
transform 1 0 93744 0 1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_833
timestamp 1669390400
transform 1 0 94640 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_96_863
timestamp 1669390400
transform 1 0 98000 0 1 78400
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_96_865
timestamp 1669390400
transform 1 0 98224 0 1 78400
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_2
timestamp 1669390400
transform 1 0 1568 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_66
timestamp 1669390400
transform 1 0 8736 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_70
timestamp 1669390400
transform 1 0 9184 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_73
timestamp 1669390400
transform 1 0 9520 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_137
timestamp 1669390400
transform 1 0 16688 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_141
timestamp 1669390400
transform 1 0 17136 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_144
timestamp 1669390400
transform 1 0 17472 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_208
timestamp 1669390400
transform 1 0 24640 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_212
timestamp 1669390400
transform 1 0 25088 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_215
timestamp 1669390400
transform 1 0 25424 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_279
timestamp 1669390400
transform 1 0 32592 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_283
timestamp 1669390400
transform 1 0 33040 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_286
timestamp 1669390400
transform 1 0 33376 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_350
timestamp 1669390400
transform 1 0 40544 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_354
timestamp 1669390400
transform 1 0 40992 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_97_357
timestamp 1669390400
transform 1 0 41328 0 -1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_421
timestamp 1669390400
transform 1 0 48496 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_425
timestamp 1669390400
transform 1 0 48944 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_428
timestamp 1669390400
transform 1 0 49280 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_458
timestamp 1669390400
transform 1 0 52640 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_465
timestamp 1669390400
transform 1 0 53424 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_469
timestamp 1669390400
transform 1 0 53872 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_478
timestamp 1669390400
transform 1 0 54880 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_485
timestamp 1669390400
transform 1 0 55664 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_489
timestamp 1669390400
transform 1 0 56112 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_493
timestamp 1669390400
transform 1 0 56560 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_496
timestamp 1669390400
transform 1 0 56896 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_499
timestamp 1669390400
transform 1 0 57232 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_532
timestamp 1669390400
transform 1 0 60928 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_536
timestamp 1669390400
transform 1 0 61376 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_540
timestamp 1669390400
transform 1 0 61824 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_559
timestamp 1669390400
transform 1 0 63952 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_563
timestamp 1669390400
transform 1 0 64400 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_567
timestamp 1669390400
transform 1 0 64848 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_97_570
timestamp 1669390400
transform 1 0 65184 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_578
timestamp 1669390400
transform 1 0 66080 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_612
timestamp 1669390400
transform 1 0 69888 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_622
timestamp 1669390400
transform 1 0 71008 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_630
timestamp 1669390400
transform 1 0 71904 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_638
timestamp 1669390400
transform 1 0 72800 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_641
timestamp 1669390400
transform 1 0 73136 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_671
timestamp 1669390400
transform 1 0 76496 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_675
timestamp 1669390400
transform 1 0 76944 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_97_679
timestamp 1669390400
transform 1 0 77392 0 -1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_97_695
timestamp 1669390400
transform 1 0 79184 0 -1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_703
timestamp 1669390400
transform 1 0 80080 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_709
timestamp 1669390400
transform 1 0 80752 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_712
timestamp 1669390400
transform 1 0 81088 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_742
timestamp 1669390400
transform 1 0 84448 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_746
timestamp 1669390400
transform 1 0 84896 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_780
timestamp 1669390400
transform 1 0 88704 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_783
timestamp 1669390400
transform 1 0 89040 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_786
timestamp 1669390400
transform 1 0 89376 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_790
timestamp 1669390400
transform 1 0 89824 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_823
timestamp 1669390400
transform 1 0 93520 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_97_840
timestamp 1669390400
transform 1 0 95424 0 -1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_848
timestamp 1669390400
transform 1 0 96320 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_854
timestamp 1669390400
transform 1 0 96992 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_97_861
timestamp 1669390400
transform 1 0 97776 0 -1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_97_865
timestamp 1669390400
transform 1 0 98224 0 -1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_98_2
timestamp 1669390400
transform 1 0 1568 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_34
timestamp 1669390400
transform 1 0 5152 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_37
timestamp 1669390400
transform 1 0 5488 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_101
timestamp 1669390400
transform 1 0 12656 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_105
timestamp 1669390400
transform 1 0 13104 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_108
timestamp 1669390400
transform 1 0 13440 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_172
timestamp 1669390400
transform 1 0 20608 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_176
timestamp 1669390400
transform 1 0 21056 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_179
timestamp 1669390400
transform 1 0 21392 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_243
timestamp 1669390400
transform 1 0 28560 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_247
timestamp 1669390400
transform 1 0 29008 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_250
timestamp 1669390400
transform 1 0 29344 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_314
timestamp 1669390400
transform 1 0 36512 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_318
timestamp 1669390400
transform 1 0 36960 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_98_321
timestamp 1669390400
transform 1 0 37296 0 1 79968
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_385
timestamp 1669390400
transform 1 0 44464 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_389
timestamp 1669390400
transform 1 0 44912 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_98_392
timestamp 1669390400
transform 1 0 45248 0 1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_424
timestamp 1669390400
transform 1 0 48832 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_457
timestamp 1669390400
transform 1 0 52528 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_463
timestamp 1669390400
transform 1 0 53200 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_493
timestamp 1669390400
transform 1 0 56560 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_500
timestamp 1669390400
transform 1 0 57344 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_98_504
timestamp 1669390400
transform 1 0 57792 0 1 79968
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_98_520
timestamp 1669390400
transform 1 0 59584 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_528
timestamp 1669390400
transform 1 0 60480 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_534
timestamp 1669390400
transform 1 0 61152 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_564
timestamp 1669390400
transform 1 0 64512 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_568
timestamp 1669390400
transform 1 0 64960 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_572
timestamp 1669390400
transform 1 0 65408 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_602
timestamp 1669390400
transform 1 0 68768 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_605
timestamp 1669390400
transform 1 0 69104 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_611
timestamp 1669390400
transform 1 0 69776 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_618
timestamp 1669390400
transform 1 0 70560 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_622
timestamp 1669390400
transform 1 0 71008 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_655
timestamp 1669390400
transform 1 0 74704 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_662
timestamp 1669390400
transform 1 0 75488 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_666
timestamp 1669390400
transform 1 0 75936 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_670
timestamp 1669390400
transform 1 0 76384 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_98_676
timestamp 1669390400
transform 1 0 77056 0 1 79968
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_684
timestamp 1669390400
transform 1 0 77952 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_688
timestamp 1669390400
transform 1 0 78400 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_719
timestamp 1669390400
transform 1 0 81872 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_723
timestamp 1669390400
transform 1 0 82320 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_730
timestamp 1669390400
transform 1 0 83104 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_737
timestamp 1669390400
transform 1 0 83888 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_744
timestamp 1669390400
transform 1 0 84672 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_747
timestamp 1669390400
transform 1 0 85008 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_750
timestamp 1669390400
transform 1 0 85344 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_754
timestamp 1669390400
transform 1 0 85792 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_758
timestamp 1669390400
transform 1 0 86240 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_762
timestamp 1669390400
transform 1 0 86688 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_764
timestamp 1669390400
transform 1 0 86912 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_815
timestamp 1669390400
transform 1 0 92624 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_818
timestamp 1669390400
transform 1 0 92960 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_821
timestamp 1669390400
transform 1 0 93296 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_98_825
timestamp 1669390400
transform 1 0 93744 0 1 79968
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_829
timestamp 1669390400
transform 1 0 94192 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_832
timestamp 1669390400
transform 1 0 94528 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_98_863
timestamp 1669390400
transform 1 0 98000 0 1 79968
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_98_865
timestamp 1669390400
transform 1 0 98224 0 1 79968
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_2
timestamp 1669390400
transform 1 0 1568 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_66
timestamp 1669390400
transform 1 0 8736 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_70
timestamp 1669390400
transform 1 0 9184 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_73
timestamp 1669390400
transform 1 0 9520 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_137
timestamp 1669390400
transform 1 0 16688 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_141
timestamp 1669390400
transform 1 0 17136 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_144
timestamp 1669390400
transform 1 0 17472 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_208
timestamp 1669390400
transform 1 0 24640 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_212
timestamp 1669390400
transform 1 0 25088 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_215
timestamp 1669390400
transform 1 0 25424 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_279
timestamp 1669390400
transform 1 0 32592 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_283
timestamp 1669390400
transform 1 0 33040 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_286
timestamp 1669390400
transform 1 0 33376 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_350
timestamp 1669390400
transform 1 0 40544 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_354
timestamp 1669390400
transform 1 0 40992 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_99_357
timestamp 1669390400
transform 1 0 41328 0 -1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_421
timestamp 1669390400
transform 1 0 48496 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_425
timestamp 1669390400
transform 1 0 48944 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_428
timestamp 1669390400
transform 1 0 49280 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_432
timestamp 1669390400
transform 1 0 49728 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_439
timestamp 1669390400
transform 1 0 50512 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_446
timestamp 1669390400
transform 1 0 51296 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_477
timestamp 1669390400
transform 1 0 54768 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_484
timestamp 1669390400
transform 1 0 55552 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_491
timestamp 1669390400
transform 1 0 56336 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_495
timestamp 1669390400
transform 1 0 56784 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_499
timestamp 1669390400
transform 1 0 57232 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_99_502
timestamp 1669390400
transform 1 0 57568 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_99_518
timestamp 1669390400
transform 1 0 59360 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_526
timestamp 1669390400
transform 1 0 60256 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_556
timestamp 1669390400
transform 1 0 63616 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_564
timestamp 1669390400
transform 1 0 64512 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_99_570
timestamp 1669390400
transform 1 0 65184 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_578
timestamp 1669390400
transform 1 0 66080 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_608
timestamp 1669390400
transform 1 0 69440 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_612
timestamp 1669390400
transform 1 0 69888 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_616
timestamp 1669390400
transform 1 0 70336 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_620
timestamp 1669390400
transform 1 0 70784 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_624
timestamp 1669390400
transform 1 0 71232 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_628
timestamp 1669390400
transform 1 0 71680 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_632
timestamp 1669390400
transform 1 0 72128 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_638
timestamp 1669390400
transform 1 0 72800 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_641
timestamp 1669390400
transform 1 0 73136 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_649
timestamp 1669390400
transform 1 0 74032 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_656
timestamp 1669390400
transform 1 0 74816 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_99_660
timestamp 1669390400
transform 1 0 75264 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_99_692
timestamp 1669390400
transform 1 0 78848 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_700
timestamp 1669390400
transform 1 0 79744 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_702
timestamp 1669390400
transform 1 0 79968 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_705
timestamp 1669390400
transform 1 0 80304 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_709
timestamp 1669390400
transform 1 0 80752 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_712
timestamp 1669390400
transform 1 0 81088 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_718
timestamp 1669390400
transform 1 0 81760 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_720
timestamp 1669390400
transform 1 0 81984 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_726
timestamp 1669390400
transform 1 0 82656 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_733
timestamp 1669390400
transform 1 0 83440 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_737
timestamp 1669390400
transform 1 0 83888 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_741
timestamp 1669390400
transform 1 0 84336 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_745
timestamp 1669390400
transform 1 0 84784 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_747
timestamp 1669390400
transform 1 0 85008 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_780
timestamp 1669390400
transform 1 0 88704 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_99_783
timestamp 1669390400
transform 1 0 89040 0 -1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_99_799
timestamp 1669390400
transform 1 0 90832 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_99_807
timestamp 1669390400
transform 1 0 91728 0 -1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_813
timestamp 1669390400
transform 1 0 92400 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_830
timestamp 1669390400
transform 1 0 94304 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_99_834
timestamp 1669390400
transform 1 0 94752 0 -1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_851
timestamp 1669390400
transform 1 0 96656 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_854
timestamp 1669390400
transform 1 0 96992 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_99_857
timestamp 1669390400
transform 1 0 97328 0 -1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_99_865
timestamp 1669390400
transform 1 0 98224 0 -1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_100_2
timestamp 1669390400
transform 1 0 1568 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_34
timestamp 1669390400
transform 1 0 5152 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_37
timestamp 1669390400
transform 1 0 5488 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_101
timestamp 1669390400
transform 1 0 12656 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_105
timestamp 1669390400
transform 1 0 13104 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_108
timestamp 1669390400
transform 1 0 13440 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_172
timestamp 1669390400
transform 1 0 20608 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_176
timestamp 1669390400
transform 1 0 21056 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_179
timestamp 1669390400
transform 1 0 21392 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_243
timestamp 1669390400
transform 1 0 28560 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_247
timestamp 1669390400
transform 1 0 29008 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_250
timestamp 1669390400
transform 1 0 29344 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_314
timestamp 1669390400
transform 1 0 36512 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_318
timestamp 1669390400
transform 1 0 36960 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_100_321
timestamp 1669390400
transform 1 0 37296 0 1 81536
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_385
timestamp 1669390400
transform 1 0 44464 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_389
timestamp 1669390400
transform 1 0 44912 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_100_392
timestamp 1669390400
transform 1 0 45248 0 1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_424
timestamp 1669390400
transform 1 0 48832 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_428
timestamp 1669390400
transform 1 0 49280 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_430
timestamp 1669390400
transform 1 0 49504 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_460
timestamp 1669390400
transform 1 0 52864 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_463
timestamp 1669390400
transform 1 0 53200 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_466
timestamp 1669390400
transform 1 0 53536 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_499
timestamp 1669390400
transform 1 0 57232 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_507
timestamp 1669390400
transform 1 0 58128 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_524
timestamp 1669390400
transform 1 0 60032 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_528
timestamp 1669390400
transform 1 0 60480 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_534
timestamp 1669390400
transform 1 0 61152 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_557
timestamp 1669390400
transform 1 0 63728 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_561
timestamp 1669390400
transform 1 0 64176 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_100_565
timestamp 1669390400
transform 1 0 64624 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_581
timestamp 1669390400
transform 1 0 66416 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_589
timestamp 1669390400
transform 1 0 67312 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_593
timestamp 1669390400
transform 1 0 67760 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_599
timestamp 1669390400
transform 1 0 68432 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_605
timestamp 1669390400
transform 1 0 69104 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_609
timestamp 1669390400
transform 1 0 69552 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_613
timestamp 1669390400
transform 1 0 70000 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_100_617
timestamp 1669390400
transform 1 0 70448 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_633
timestamp 1669390400
transform 1 0 72240 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_645
timestamp 1669390400
transform 1 0 73584 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_649
timestamp 1669390400
transform 1 0 74032 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_653
timestamp 1669390400
transform 1 0 74480 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_663
timestamp 1669390400
transform 1 0 75600 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_673
timestamp 1669390400
transform 1 0 76720 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_676
timestamp 1669390400
transform 1 0 77056 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_100_685
timestamp 1669390400
transform 1 0 78064 0 1 81536
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_701
timestamp 1669390400
transform 1 0 79856 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_705
timestamp 1669390400
transform 1 0 80304 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_707
timestamp 1669390400
transform 1 0 80528 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_710
timestamp 1669390400
transform 1 0 80864 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_717
timestamp 1669390400
transform 1 0 81648 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_100_721
timestamp 1669390400
transform 1 0 82096 0 1 81536
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_725
timestamp 1669390400
transform 1 0 82544 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_731
timestamp 1669390400
transform 1 0 83216 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_738
timestamp 1669390400
transform 1 0 84000 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_742
timestamp 1669390400
transform 1 0 84448 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_744
timestamp 1669390400
transform 1 0 84672 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_747
timestamp 1669390400
transform 1 0 85008 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_798
timestamp 1669390400
transform 1 0 90720 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_100_802
timestamp 1669390400
transform 1 0 91168 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_810
timestamp 1669390400
transform 1 0 92064 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_812
timestamp 1669390400
transform 1 0 92288 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_815
timestamp 1669390400
transform 1 0 92624 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_818
timestamp 1669390400
transform 1 0 92960 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_834
timestamp 1669390400
transform 1 0 94752 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_851
timestamp 1669390400
transform 1 0 96656 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_855
timestamp 1669390400
transform 1 0 97104 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_859
timestamp 1669390400
transform 1 0 97552 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_100_863
timestamp 1669390400
transform 1 0 98000 0 1 81536
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_100_865
timestamp 1669390400
transform 1 0 98224 0 1 81536
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_2
timestamp 1669390400
transform 1 0 1568 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_66
timestamp 1669390400
transform 1 0 8736 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_70
timestamp 1669390400
transform 1 0 9184 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_73
timestamp 1669390400
transform 1 0 9520 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_137
timestamp 1669390400
transform 1 0 16688 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_141
timestamp 1669390400
transform 1 0 17136 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_144
timestamp 1669390400
transform 1 0 17472 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_208
timestamp 1669390400
transform 1 0 24640 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_212
timestamp 1669390400
transform 1 0 25088 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_215
timestamp 1669390400
transform 1 0 25424 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_279
timestamp 1669390400
transform 1 0 32592 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_283
timestamp 1669390400
transform 1 0 33040 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_286
timestamp 1669390400
transform 1 0 33376 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_350
timestamp 1669390400
transform 1 0 40544 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_354
timestamp 1669390400
transform 1 0 40992 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_101_357
timestamp 1669390400
transform 1 0 41328 0 -1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_421
timestamp 1669390400
transform 1 0 48496 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_425
timestamp 1669390400
transform 1 0 48944 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_101_428
timestamp 1669390400
transform 1 0 49280 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_444
timestamp 1669390400
transform 1 0 51072 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_496
timestamp 1669390400
transform 1 0 56896 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_499
timestamp 1669390400
transform 1 0 57232 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_529
timestamp 1669390400
transform 1 0 60592 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_533
timestamp 1669390400
transform 1 0 61040 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_543
timestamp 1669390400
transform 1 0 62160 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_551
timestamp 1669390400
transform 1 0 63056 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_559
timestamp 1669390400
transform 1 0 63952 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_567
timestamp 1669390400
transform 1 0 64848 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_101_570
timestamp 1669390400
transform 1 0 65184 0 -1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_602
timestamp 1669390400
transform 1 0 68768 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_606
timestamp 1669390400
transform 1 0 69216 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_610
timestamp 1669390400
transform 1 0 69664 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_101_614
timestamp 1669390400
transform 1 0 70112 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_630
timestamp 1669390400
transform 1 0 71904 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_638
timestamp 1669390400
transform 1 0 72800 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_641
timestamp 1669390400
transform 1 0 73136 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_645
timestamp 1669390400
transform 1 0 73584 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_649
timestamp 1669390400
transform 1 0 74032 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_653
timestamp 1669390400
transform 1 0 74480 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_655
timestamp 1669390400
transform 1 0 74704 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_658
timestamp 1669390400
transform 1 0 75040 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_689
timestamp 1669390400
transform 1 0 78512 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_693
timestamp 1669390400
transform 1 0 78960 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_701
timestamp 1669390400
transform 1 0 79856 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_703
timestamp 1669390400
transform 1 0 80080 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_709
timestamp 1669390400
transform 1 0 80752 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_712
timestamp 1669390400
transform 1 0 81088 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_716
timestamp 1669390400
transform 1 0 81536 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_747
timestamp 1669390400
transform 1 0 85008 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_751
timestamp 1669390400
transform 1 0 85456 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_755
timestamp 1669390400
transform 1 0 85904 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_759
timestamp 1669390400
transform 1 0 86352 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_101_763
timestamp 1669390400
transform 1 0 86800 0 -1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_779
timestamp 1669390400
transform 1 0 88592 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_783
timestamp 1669390400
transform 1 0 89040 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_791
timestamp 1669390400
transform 1 0 89936 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_795
timestamp 1669390400
transform 1 0 90384 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_101_799
timestamp 1669390400
transform 1 0 90832 0 -1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_101_851
timestamp 1669390400
transform 1 0 96656 0 -1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_101_854
timestamp 1669390400
transform 1 0 96992 0 -1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_101_862
timestamp 1669390400
transform 1 0 97888 0 -1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_102_2
timestamp 1669390400
transform 1 0 1568 0 1 83104
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_34
timestamp 1669390400
transform 1 0 5152 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_37
timestamp 1669390400
transform 1 0 5488 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_101
timestamp 1669390400
transform 1 0 12656 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_105
timestamp 1669390400
transform 1 0 13104 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_108
timestamp 1669390400
transform 1 0 13440 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_172
timestamp 1669390400
transform 1 0 20608 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_176
timestamp 1669390400
transform 1 0 21056 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_179
timestamp 1669390400
transform 1 0 21392 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_243
timestamp 1669390400
transform 1 0 28560 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_247
timestamp 1669390400
transform 1 0 29008 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_250
timestamp 1669390400
transform 1 0 29344 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_314
timestamp 1669390400
transform 1 0 36512 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_318
timestamp 1669390400
transform 1 0 36960 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_321
timestamp 1669390400
transform 1 0 37296 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_385
timestamp 1669390400
transform 1 0 44464 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_389
timestamp 1669390400
transform 1 0 44912 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_102_392
timestamp 1669390400
transform 1 0 45248 0 1 83104
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_456
timestamp 1669390400
transform 1 0 52416 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_460
timestamp 1669390400
transform 1 0 52864 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_463
timestamp 1669390400
transform 1 0 53200 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_469
timestamp 1669390400
transform 1 0 53872 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_476
timestamp 1669390400
transform 1 0 54656 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_480
timestamp 1669390400
transform 1 0 55104 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_498
timestamp 1669390400
transform 1 0 57120 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_502
timestamp 1669390400
transform 1 0 57568 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_509
timestamp 1669390400
transform 1 0 58352 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_525
timestamp 1669390400
transform 1 0 60144 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_529
timestamp 1669390400
transform 1 0 60592 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_531
timestamp 1669390400
transform 1 0 60816 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_534
timestamp 1669390400
transform 1 0 61152 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_550
timestamp 1669390400
transform 1 0 62944 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_567
timestamp 1669390400
transform 1 0 64848 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_571
timestamp 1669390400
transform 1 0 65296 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_587
timestamp 1669390400
transform 1 0 67088 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_591
timestamp 1669390400
transform 1 0 67536 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_102_594
timestamp 1669390400
transform 1 0 67872 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_602
timestamp 1669390400
transform 1 0 68768 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_605
timestamp 1669390400
transform 1 0 69104 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_612
timestamp 1669390400
transform 1 0 69888 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_620
timestamp 1669390400
transform 1 0 70784 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_624
timestamp 1669390400
transform 1 0 71232 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_626
timestamp 1669390400
transform 1 0 71456 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_629
timestamp 1669390400
transform 1 0 71792 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_633
timestamp 1669390400
transform 1 0 72240 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_643
timestamp 1669390400
transform 1 0 73360 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_647
timestamp 1669390400
transform 1 0 73808 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_664
timestamp 1669390400
transform 1 0 75712 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_672
timestamp 1669390400
transform 1 0 76608 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_676
timestamp 1669390400
transform 1 0 77056 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_692
timestamp 1669390400
transform 1 0 78848 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_696
timestamp 1669390400
transform 1 0 79296 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_700
timestamp 1669390400
transform 1 0 79744 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_731
timestamp 1669390400
transform 1 0 83216 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_738
timestamp 1669390400
transform 1 0 84000 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_742
timestamp 1669390400
transform 1 0 84448 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_744
timestamp 1669390400
transform 1 0 84672 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_747
timestamp 1669390400
transform 1 0 85008 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_750
timestamp 1669390400
transform 1 0 85344 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_102_754
timestamp 1669390400
transform 1 0 85792 0 1 83104
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_772
timestamp 1669390400
transform 1 0 87808 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_789
timestamp 1669390400
transform 1 0 89712 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_793
timestamp 1669390400
transform 1 0 90160 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_795
timestamp 1669390400
transform 1 0 90384 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_798
timestamp 1669390400
transform 1 0 90720 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_815
timestamp 1669390400
transform 1 0 92624 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_818
timestamp 1669390400
transform 1 0 92960 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_102_825
timestamp 1669390400
transform 1 0 93744 0 1 83104
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_829
timestamp 1669390400
transform 1 0 94192 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_832
timestamp 1669390400
transform 1 0 94528 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_102_863
timestamp 1669390400
transform 1 0 98000 0 1 83104
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_102_865
timestamp 1669390400
transform 1 0 98224 0 1 83104
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_2
timestamp 1669390400
transform 1 0 1568 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_66
timestamp 1669390400
transform 1 0 8736 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_70
timestamp 1669390400
transform 1 0 9184 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_73
timestamp 1669390400
transform 1 0 9520 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_137
timestamp 1669390400
transform 1 0 16688 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_141
timestamp 1669390400
transform 1 0 17136 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_144
timestamp 1669390400
transform 1 0 17472 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_208
timestamp 1669390400
transform 1 0 24640 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_212
timestamp 1669390400
transform 1 0 25088 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_215
timestamp 1669390400
transform 1 0 25424 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_279
timestamp 1669390400
transform 1 0 32592 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_283
timestamp 1669390400
transform 1 0 33040 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_286
timestamp 1669390400
transform 1 0 33376 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_350
timestamp 1669390400
transform 1 0 40544 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_354
timestamp 1669390400
transform 1 0 40992 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_103_357
timestamp 1669390400
transform 1 0 41328 0 -1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_421
timestamp 1669390400
transform 1 0 48496 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_425
timestamp 1669390400
transform 1 0 48944 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_103_428
timestamp 1669390400
transform 1 0 49280 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_436
timestamp 1669390400
transform 1 0 50176 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_440
timestamp 1669390400
transform 1 0 50624 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_471
timestamp 1669390400
transform 1 0 54096 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_475
timestamp 1669390400
transform 1 0 54544 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_103_479
timestamp 1669390400
transform 1 0 54992 0 -1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_495
timestamp 1669390400
transform 1 0 56784 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_499
timestamp 1669390400
transform 1 0 57232 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_103_502
timestamp 1669390400
transform 1 0 57568 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_560
timestamp 1669390400
transform 1 0 64064 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_564
timestamp 1669390400
transform 1 0 64512 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_570
timestamp 1669390400
transform 1 0 65184 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_574
timestamp 1669390400
transform 1 0 65632 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_577
timestamp 1669390400
transform 1 0 65968 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_608
timestamp 1669390400
transform 1 0 69440 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_627
timestamp 1669390400
transform 1 0 71568 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_637
timestamp 1669390400
transform 1 0 72688 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_641
timestamp 1669390400
transform 1 0 73136 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_672
timestamp 1669390400
transform 1 0 76608 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_676
timestamp 1669390400
transform 1 0 77056 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_706
timestamp 1669390400
transform 1 0 80416 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_712
timestamp 1669390400
transform 1 0 81088 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_742
timestamp 1669390400
transform 1 0 84448 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_749
timestamp 1669390400
transform 1 0 85232 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_780
timestamp 1669390400
transform 1 0 88704 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_783
timestamp 1669390400
transform 1 0 89040 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_790
timestamp 1669390400
transform 1 0 89824 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_794
timestamp 1669390400
transform 1 0 90272 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_798
timestamp 1669390400
transform 1 0 90720 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_802
timestamp 1669390400
transform 1 0 91168 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_103_833
timestamp 1669390400
transform 1 0 94640 0 -1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_835
timestamp 1669390400
transform 1 0 94864 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_103_851
timestamp 1669390400
transform 1 0 96656 0 -1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_103_854
timestamp 1669390400
transform 1 0 96992 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_103_862
timestamp 1669390400
transform 1 0 97888 0 -1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_2
timestamp 1669390400
transform 1 0 1568 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_34
timestamp 1669390400
transform 1 0 5152 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_37
timestamp 1669390400
transform 1 0 5488 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_101
timestamp 1669390400
transform 1 0 12656 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_105
timestamp 1669390400
transform 1 0 13104 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_108
timestamp 1669390400
transform 1 0 13440 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_172
timestamp 1669390400
transform 1 0 20608 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_176
timestamp 1669390400
transform 1 0 21056 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_179
timestamp 1669390400
transform 1 0 21392 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_243
timestamp 1669390400
transform 1 0 28560 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_247
timestamp 1669390400
transform 1 0 29008 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_250
timestamp 1669390400
transform 1 0 29344 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_314
timestamp 1669390400
transform 1 0 36512 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_318
timestamp 1669390400
transform 1 0 36960 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_104_321
timestamp 1669390400
transform 1 0 37296 0 1 84672
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_385
timestamp 1669390400
transform 1 0 44464 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_389
timestamp 1669390400
transform 1 0 44912 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_104_392
timestamp 1669390400
transform 1 0 45248 0 1 84672
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_104_424
timestamp 1669390400
transform 1 0 48832 0 1 84672
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_440
timestamp 1669390400
transform 1 0 50624 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_448
timestamp 1669390400
transform 1 0 51520 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_452
timestamp 1669390400
transform 1 0 51968 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_459
timestamp 1669390400
transform 1 0 52752 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_463
timestamp 1669390400
transform 1 0 53200 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_467
timestamp 1669390400
transform 1 0 53648 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_470
timestamp 1669390400
transform 1 0 53984 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_501
timestamp 1669390400
transform 1 0 57456 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_505
timestamp 1669390400
transform 1 0 57904 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_524
timestamp 1669390400
transform 1 0 60032 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_528
timestamp 1669390400
transform 1 0 60480 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_534
timestamp 1669390400
transform 1 0 61152 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_541
timestamp 1669390400
transform 1 0 61936 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_545
timestamp 1669390400
transform 1 0 62384 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_575
timestamp 1669390400
transform 1 0 65744 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_592
timestamp 1669390400
transform 1 0 67648 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_600
timestamp 1669390400
transform 1 0 68544 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_602
timestamp 1669390400
transform 1 0 68768 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_605
timestamp 1669390400
transform 1 0 69104 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_635
timestamp 1669390400
transform 1 0 72464 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_639
timestamp 1669390400
transform 1 0 72912 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_643
timestamp 1669390400
transform 1 0 73360 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_653
timestamp 1669390400
transform 1 0 74480 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_670
timestamp 1669390400
transform 1 0 76384 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_676
timestamp 1669390400
transform 1 0 77056 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_727
timestamp 1669390400
transform 1 0 82768 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_731
timestamp 1669390400
transform 1 0 83216 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_104_735
timestamp 1669390400
transform 1 0 83664 0 1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_743
timestamp 1669390400
transform 1 0 84560 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_747
timestamp 1669390400
transform 1 0 85008 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_777
timestamp 1669390400
transform 1 0 88368 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_794
timestamp 1669390400
transform 1 0 90272 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_798
timestamp 1669390400
transform 1 0 90720 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_815
timestamp 1669390400
transform 1 0 92624 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_818
timestamp 1669390400
transform 1 0 92960 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_104_825
timestamp 1669390400
transform 1 0 93744 0 1 84672
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_829
timestamp 1669390400
transform 1 0 94192 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_832
timestamp 1669390400
transform 1 0 94528 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_104_863
timestamp 1669390400
transform 1 0 98000 0 1 84672
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_104_865
timestamp 1669390400
transform 1 0 98224 0 1 84672
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_2
timestamp 1669390400
transform 1 0 1568 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_66
timestamp 1669390400
transform 1 0 8736 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_70
timestamp 1669390400
transform 1 0 9184 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_73
timestamp 1669390400
transform 1 0 9520 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_137
timestamp 1669390400
transform 1 0 16688 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_141
timestamp 1669390400
transform 1 0 17136 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_144
timestamp 1669390400
transform 1 0 17472 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_208
timestamp 1669390400
transform 1 0 24640 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_212
timestamp 1669390400
transform 1 0 25088 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_215
timestamp 1669390400
transform 1 0 25424 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_279
timestamp 1669390400
transform 1 0 32592 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_283
timestamp 1669390400
transform 1 0 33040 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_286
timestamp 1669390400
transform 1 0 33376 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_350
timestamp 1669390400
transform 1 0 40544 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_354
timestamp 1669390400
transform 1 0 40992 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_105_357
timestamp 1669390400
transform 1 0 41328 0 -1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_421
timestamp 1669390400
transform 1 0 48496 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_425
timestamp 1669390400
transform 1 0 48944 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_105_428
timestamp 1669390400
transform 1 0 49280 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_436
timestamp 1669390400
transform 1 0 50176 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_440
timestamp 1669390400
transform 1 0 50624 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_442
timestamp 1669390400
transform 1 0 50848 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_472
timestamp 1669390400
transform 1 0 54208 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_476
timestamp 1669390400
transform 1 0 54656 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_480
timestamp 1669390400
transform 1 0 55104 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_496
timestamp 1669390400
transform 1 0 56896 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_499
timestamp 1669390400
transform 1 0 57232 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_529
timestamp 1669390400
transform 1 0 60592 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_560
timestamp 1669390400
transform 1 0 64064 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_564
timestamp 1669390400
transform 1 0 64512 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_570
timestamp 1669390400
transform 1 0 65184 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_574
timestamp 1669390400
transform 1 0 65632 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_626
timestamp 1669390400
transform 1 0 71456 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_630
timestamp 1669390400
transform 1 0 71904 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_634
timestamp 1669390400
transform 1 0 72352 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_638
timestamp 1669390400
transform 1 0 72800 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_641
timestamp 1669390400
transform 1 0 73136 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_650
timestamp 1669390400
transform 1 0 74144 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_681
timestamp 1669390400
transform 1 0 77616 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_698
timestamp 1669390400
transform 1 0 79520 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_702
timestamp 1669390400
transform 1 0 79968 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_708
timestamp 1669390400
transform 1 0 80640 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_712
timestamp 1669390400
transform 1 0 81088 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_742
timestamp 1669390400
transform 1 0 84448 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_746
timestamp 1669390400
transform 1 0 84896 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_750
timestamp 1669390400
transform 1 0 85344 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_780
timestamp 1669390400
transform 1 0 88704 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_783
timestamp 1669390400
transform 1 0 89040 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_105_786
timestamp 1669390400
transform 1 0 89376 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_794
timestamp 1669390400
transform 1 0 90272 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_105_825
timestamp 1669390400
transform 1 0 93744 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_833
timestamp 1669390400
transform 1 0 94640 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_837
timestamp 1669390400
transform 1 0 95088 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_105_839
timestamp 1669390400
transform 1 0 95312 0 -1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_846
timestamp 1669390400
transform 1 0 96096 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_105_850
timestamp 1669390400
transform 1 0 96544 0 -1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_105_854
timestamp 1669390400
transform 1 0 96992 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_105_862
timestamp 1669390400
transform 1 0 97888 0 -1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_2
timestamp 1669390400
transform 1 0 1568 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_34
timestamp 1669390400
transform 1 0 5152 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_37
timestamp 1669390400
transform 1 0 5488 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_101
timestamp 1669390400
transform 1 0 12656 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_105
timestamp 1669390400
transform 1 0 13104 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_108
timestamp 1669390400
transform 1 0 13440 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_172
timestamp 1669390400
transform 1 0 20608 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_176
timestamp 1669390400
transform 1 0 21056 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_179
timestamp 1669390400
transform 1 0 21392 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_243
timestamp 1669390400
transform 1 0 28560 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_247
timestamp 1669390400
transform 1 0 29008 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_250
timestamp 1669390400
transform 1 0 29344 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_314
timestamp 1669390400
transform 1 0 36512 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_318
timestamp 1669390400
transform 1 0 36960 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_106_321
timestamp 1669390400
transform 1 0 37296 0 1 86240
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_385
timestamp 1669390400
transform 1 0 44464 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_389
timestamp 1669390400
transform 1 0 44912 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_106_392
timestamp 1669390400
transform 1 0 45248 0 1 86240
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_424
timestamp 1669390400
transform 1 0 48832 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_440
timestamp 1669390400
transform 1 0 50624 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_448
timestamp 1669390400
transform 1 0 51520 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_452
timestamp 1669390400
transform 1 0 51968 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_459
timestamp 1669390400
transform 1 0 52752 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_463
timestamp 1669390400
transform 1 0 53200 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_479
timestamp 1669390400
transform 1 0 54992 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_487
timestamp 1669390400
transform 1 0 55888 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_489
timestamp 1669390400
transform 1 0 56112 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_519
timestamp 1669390400
transform 1 0 59472 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_527
timestamp 1669390400
transform 1 0 60368 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_531
timestamp 1669390400
transform 1 0 60816 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_534
timestamp 1669390400
transform 1 0 61152 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_541
timestamp 1669390400
transform 1 0 61936 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_545
timestamp 1669390400
transform 1 0 62384 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_547
timestamp 1669390400
transform 1 0 62608 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_577
timestamp 1669390400
transform 1 0 65968 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_581
timestamp 1669390400
transform 1 0 66416 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_585
timestamp 1669390400
transform 1 0 66864 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_593
timestamp 1669390400
transform 1 0 67760 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_595
timestamp 1669390400
transform 1 0 67984 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_602
timestamp 1669390400
transform 1 0 68768 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_605
timestamp 1669390400
transform 1 0 69104 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_621
timestamp 1669390400
transform 1 0 70896 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_638
timestamp 1669390400
transform 1 0 72800 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_648
timestamp 1669390400
transform 1 0 73920 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_658
timestamp 1669390400
transform 1 0 75040 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_666
timestamp 1669390400
transform 1 0 75936 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_672
timestamp 1669390400
transform 1 0 76608 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_676
timestamp 1669390400
transform 1 0 77056 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_679
timestamp 1669390400
transform 1 0 77392 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_687
timestamp 1669390400
transform 1 0 78288 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_691
timestamp 1669390400
transform 1 0 78736 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_695
timestamp 1669390400
transform 1 0 79184 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_697
timestamp 1669390400
transform 1 0 79408 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_700
timestamp 1669390400
transform 1 0 79744 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_708
timestamp 1669390400
transform 1 0 80640 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_714
timestamp 1669390400
transform 1 0 81312 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_721
timestamp 1669390400
transform 1 0 82096 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_728
timestamp 1669390400
transform 1 0 82880 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_732
timestamp 1669390400
transform 1 0 83328 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_740
timestamp 1669390400
transform 1 0 84224 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_744
timestamp 1669390400
transform 1 0 84672 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_106_747
timestamp 1669390400
transform 1 0 85008 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_755
timestamp 1669390400
transform 1 0 85904 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_762
timestamp 1669390400
transform 1 0 86688 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_766
timestamp 1669390400
transform 1 0 87136 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_783
timestamp 1669390400
transform 1 0 89040 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_787
timestamp 1669390400
transform 1 0 89488 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_106_803
timestamp 1669390400
transform 1 0 91280 0 1 86240
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_810
timestamp 1669390400
transform 1 0 92064 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_814
timestamp 1669390400
transform 1 0 92512 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_818
timestamp 1669390400
transform 1 0 92960 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_834
timestamp 1669390400
transform 1 0 94752 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_106_838
timestamp 1669390400
transform 1 0 95200 0 1 86240
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_106_846
timestamp 1669390400
transform 1 0 96096 0 1 86240
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_106_862
timestamp 1669390400
transform 1 0 97888 0 1 86240
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_2
timestamp 1669390400
transform 1 0 1568 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_5
timestamp 1669390400
transform 1 0 1904 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_69
timestamp 1669390400
transform 1 0 9072 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_73
timestamp 1669390400
transform 1 0 9520 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_137
timestamp 1669390400
transform 1 0 16688 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_141
timestamp 1669390400
transform 1 0 17136 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_144
timestamp 1669390400
transform 1 0 17472 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_208
timestamp 1669390400
transform 1 0 24640 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_212
timestamp 1669390400
transform 1 0 25088 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_215
timestamp 1669390400
transform 1 0 25424 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_279
timestamp 1669390400
transform 1 0 32592 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_283
timestamp 1669390400
transform 1 0 33040 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_286
timestamp 1669390400
transform 1 0 33376 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_350
timestamp 1669390400
transform 1 0 40544 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_354
timestamp 1669390400
transform 1 0 40992 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_107_357
timestamp 1669390400
transform 1 0 41328 0 -1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_421
timestamp 1669390400
transform 1 0 48496 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_425
timestamp 1669390400
transform 1 0 48944 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_107_428
timestamp 1669390400
transform 1 0 49280 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_460
timestamp 1669390400
transform 1 0 52864 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_476
timestamp 1669390400
transform 1 0 54656 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_478
timestamp 1669390400
transform 1 0 54880 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_481
timestamp 1669390400
transform 1 0 55216 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_485
timestamp 1669390400
transform 1 0 55664 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_489
timestamp 1669390400
transform 1 0 56112 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_499
timestamp 1669390400
transform 1 0 57232 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_502
timestamp 1669390400
transform 1 0 57568 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_519
timestamp 1669390400
transform 1 0 59472 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_550
timestamp 1669390400
transform 1 0 62944 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_567
timestamp 1669390400
transform 1 0 64848 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_570
timestamp 1669390400
transform 1 0 65184 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_573
timestamp 1669390400
transform 1 0 65520 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_581
timestamp 1669390400
transform 1 0 66416 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_585
timestamp 1669390400
transform 1 0 66864 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_587
timestamp 1669390400
transform 1 0 67088 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_617
timestamp 1669390400
transform 1 0 70448 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_621
timestamp 1669390400
transform 1 0 70896 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_638
timestamp 1669390400
transform 1 0 72800 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_641
timestamp 1669390400
transform 1 0 73136 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_644
timestamp 1669390400
transform 1 0 73472 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_648
timestamp 1669390400
transform 1 0 73920 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_652
timestamp 1669390400
transform 1 0 74368 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_655
timestamp 1669390400
transform 1 0 74704 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_659
timestamp 1669390400
transform 1 0 75152 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_107_663
timestamp 1669390400
transform 1 0 75600 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_695
timestamp 1669390400
transform 1 0 79184 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_703
timestamp 1669390400
transform 1 0 80080 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_707
timestamp 1669390400
transform 1 0 80528 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_709
timestamp 1669390400
transform 1 0 80752 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_107_712
timestamp 1669390400
transform 1 0 81088 0 -1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_107_744
timestamp 1669390400
transform 1 0 84672 0 -1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_760
timestamp 1669390400
transform 1 0 86464 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_762
timestamp 1669390400
transform 1 0 86688 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_769
timestamp 1669390400
transform 1 0 87472 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_777
timestamp 1669390400
transform 1 0 88368 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_107_783
timestamp 1669390400
transform 1 0 89040 0 -1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_834
timestamp 1669390400
transform 1 0 94752 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_838
timestamp 1669390400
transform 1 0 95200 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_846
timestamp 1669390400
transform 1 0 96096 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_107_850
timestamp 1669390400
transform 1 0 96544 0 -1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_107_854
timestamp 1669390400
transform 1 0 96992 0 -1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_107_862
timestamp 1669390400
transform 1 0 97888 0 -1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_2
timestamp 1669390400
transform 1 0 1568 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_19
timestamp 1669390400
transform 1 0 3472 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_37
timestamp 1669390400
transform 1 0 5488 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_101
timestamp 1669390400
transform 1 0 12656 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_105
timestamp 1669390400
transform 1 0 13104 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_108
timestamp 1669390400
transform 1 0 13440 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_172
timestamp 1669390400
transform 1 0 20608 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_176
timestamp 1669390400
transform 1 0 21056 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_179
timestamp 1669390400
transform 1 0 21392 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_243
timestamp 1669390400
transform 1 0 28560 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_247
timestamp 1669390400
transform 1 0 29008 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_250
timestamp 1669390400
transform 1 0 29344 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_314
timestamp 1669390400
transform 1 0 36512 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_318
timestamp 1669390400
transform 1 0 36960 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_321
timestamp 1669390400
transform 1 0 37296 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_385
timestamp 1669390400
transform 1 0 44464 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_389
timestamp 1669390400
transform 1 0 44912 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_392
timestamp 1669390400
transform 1 0 45248 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_456
timestamp 1669390400
transform 1 0 52416 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_460
timestamp 1669390400
transform 1 0 52864 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_463
timestamp 1669390400
transform 1 0 53200 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_471
timestamp 1669390400
transform 1 0 54096 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_475
timestamp 1669390400
transform 1 0 54544 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_478
timestamp 1669390400
transform 1 0 54880 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_494
timestamp 1669390400
transform 1 0 56672 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_498
timestamp 1669390400
transform 1 0 57120 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_505
timestamp 1669390400
transform 1 0 57904 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_513
timestamp 1669390400
transform 1 0 58800 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_517
timestamp 1669390400
transform 1 0 59248 0 1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_521
timestamp 1669390400
transform 1 0 59696 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_531
timestamp 1669390400
transform 1 0 60816 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_534
timestamp 1669390400
transform 1 0 61152 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_550
timestamp 1669390400
transform 1 0 62944 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_560
timestamp 1669390400
transform 1 0 64064 0 1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_108_564
timestamp 1669390400
transform 1 0 64512 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_596
timestamp 1669390400
transform 1 0 68096 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_600
timestamp 1669390400
transform 1 0 68544 0 1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_602
timestamp 1669390400
transform 1 0 68768 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_108_605
timestamp 1669390400
transform 1 0 69104 0 1 87808
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_613
timestamp 1669390400
transform 1 0 70000 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_619
timestamp 1669390400
transform 1 0 70672 0 1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_108_623
timestamp 1669390400
transform 1 0 71120 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_655
timestamp 1669390400
transform 1 0 74704 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_108_671
timestamp 1669390400
transform 1 0 76496 0 1 87808
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_673
timestamp 1669390400
transform 1 0 76720 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_676
timestamp 1669390400
transform 1 0 77056 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_740
timestamp 1669390400
transform 1 0 84224 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_744
timestamp 1669390400
transform 1 0 84672 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_108_747
timestamp 1669390400
transform 1 0 85008 0 1 87808
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_108_811
timestamp 1669390400
transform 1 0 92176 0 1 87808
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_108_815
timestamp 1669390400
transform 1 0 92624 0 1 87808
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_108_818
timestamp 1669390400
transform 1 0 92960 0 1 87808
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_108_850
timestamp 1669390400
transform 1 0 96544 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_2
timestamp 1669390400
transform 1 0 1568 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_66
timestamp 1669390400
transform 1 0 8736 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_70
timestamp 1669390400
transform 1 0 9184 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_73
timestamp 1669390400
transform 1 0 9520 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_137
timestamp 1669390400
transform 1 0 16688 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_141
timestamp 1669390400
transform 1 0 17136 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_144
timestamp 1669390400
transform 1 0 17472 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_208
timestamp 1669390400
transform 1 0 24640 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_212
timestamp 1669390400
transform 1 0 25088 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_215
timestamp 1669390400
transform 1 0 25424 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_279
timestamp 1669390400
transform 1 0 32592 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_283
timestamp 1669390400
transform 1 0 33040 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_286
timestamp 1669390400
transform 1 0 33376 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_350
timestamp 1669390400
transform 1 0 40544 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_354
timestamp 1669390400
transform 1 0 40992 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_357
timestamp 1669390400
transform 1 0 41328 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_421
timestamp 1669390400
transform 1 0 48496 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_425
timestamp 1669390400
transform 1 0 48944 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_428
timestamp 1669390400
transform 1 0 49280 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_492
timestamp 1669390400
transform 1 0 56448 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_496
timestamp 1669390400
transform 1 0 56896 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_109_499
timestamp 1669390400
transform 1 0 57232 0 -1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_531
timestamp 1669390400
transform 1 0 60816 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_547
timestamp 1669390400
transform 1 0 62608 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_549
timestamp 1669390400
transform 1 0 62832 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_552
timestamp 1669390400
transform 1 0 63168 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_556
timestamp 1669390400
transform 1 0 63616 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_564
timestamp 1669390400
transform 1 0 64512 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_570
timestamp 1669390400
transform 1 0 65184 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_586
timestamp 1669390400
transform 1 0 66976 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_594
timestamp 1669390400
transform 1 0 67872 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_624
timestamp 1669390400
transform 1 0 71232 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_628
timestamp 1669390400
transform 1 0 71680 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_636
timestamp 1669390400
transform 1 0 72576 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_638
timestamp 1669390400
transform 1 0 72800 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_641
timestamp 1669390400
transform 1 0 73136 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_705
timestamp 1669390400
transform 1 0 80304 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_709
timestamp 1669390400
transform 1 0 80752 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_109_712
timestamp 1669390400
transform 1 0 81088 0 -1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_776
timestamp 1669390400
transform 1 0 88256 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_780
timestamp 1669390400
transform 1 0 88704 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_783
timestamp 1669390400
transform 1 0 89040 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_791
timestamp 1669390400
transform 1 0 89936 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_109_795
timestamp 1669390400
transform 1 0 90384 0 -1 89376
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_797
timestamp 1669390400
transform 1 0 90608 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_109_827
timestamp 1669390400
transform 1 0 93968 0 -1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_843
timestamp 1669390400
transform 1 0 95760 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_109_851
timestamp 1669390400
transform 1 0 96656 0 -1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_109_854
timestamp 1669390400
transform 1 0 96992 0 -1 89376
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_109_862
timestamp 1669390400
transform 1 0 97888 0 -1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_2
timestamp 1669390400
transform 1 0 1568 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_34
timestamp 1669390400
transform 1 0 5152 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_37
timestamp 1669390400
transform 1 0 5488 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_101
timestamp 1669390400
transform 1 0 12656 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_105
timestamp 1669390400
transform 1 0 13104 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_108
timestamp 1669390400
transform 1 0 13440 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_172
timestamp 1669390400
transform 1 0 20608 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_176
timestamp 1669390400
transform 1 0 21056 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_179
timestamp 1669390400
transform 1 0 21392 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_243
timestamp 1669390400
transform 1 0 28560 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_247
timestamp 1669390400
transform 1 0 29008 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_250
timestamp 1669390400
transform 1 0 29344 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_314
timestamp 1669390400
transform 1 0 36512 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_318
timestamp 1669390400
transform 1 0 36960 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_321
timestamp 1669390400
transform 1 0 37296 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_385
timestamp 1669390400
transform 1 0 44464 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_389
timestamp 1669390400
transform 1 0 44912 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_392
timestamp 1669390400
transform 1 0 45248 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_456
timestamp 1669390400
transform 1 0 52416 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_460
timestamp 1669390400
transform 1 0 52864 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_463
timestamp 1669390400
transform 1 0 53200 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_527
timestamp 1669390400
transform 1 0 60368 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_531
timestamp 1669390400
transform 1 0 60816 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_534
timestamp 1669390400
transform 1 0 61152 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_598
timestamp 1669390400
transform 1 0 68320 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_602
timestamp 1669390400
transform 1 0 68768 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_605
timestamp 1669390400
transform 1 0 69104 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_669
timestamp 1669390400
transform 1 0 76272 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_673
timestamp 1669390400
transform 1 0 76720 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_676
timestamp 1669390400
transform 1 0 77056 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_740
timestamp 1669390400
transform 1 0 84224 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_744
timestamp 1669390400
transform 1 0 84672 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_110_747
timestamp 1669390400
transform 1 0 85008 0 1 89376
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_110_811
timestamp 1669390400
transform 1 0 92176 0 1 89376
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_110_815
timestamp 1669390400
transform 1 0 92624 0 1 89376
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_110_818
timestamp 1669390400
transform 1 0 92960 0 1 89376
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_110_850
timestamp 1669390400
transform 1 0 96544 0 1 89376
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_2
timestamp 1669390400
transform 1 0 1568 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_66
timestamp 1669390400
transform 1 0 8736 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_70
timestamp 1669390400
transform 1 0 9184 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_73
timestamp 1669390400
transform 1 0 9520 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_137
timestamp 1669390400
transform 1 0 16688 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_141
timestamp 1669390400
transform 1 0 17136 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_144
timestamp 1669390400
transform 1 0 17472 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_208
timestamp 1669390400
transform 1 0 24640 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_212
timestamp 1669390400
transform 1 0 25088 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_215
timestamp 1669390400
transform 1 0 25424 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_279
timestamp 1669390400
transform 1 0 32592 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_283
timestamp 1669390400
transform 1 0 33040 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_286
timestamp 1669390400
transform 1 0 33376 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_350
timestamp 1669390400
transform 1 0 40544 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_354
timestamp 1669390400
transform 1 0 40992 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_357
timestamp 1669390400
transform 1 0 41328 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_421
timestamp 1669390400
transform 1 0 48496 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_425
timestamp 1669390400
transform 1 0 48944 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_428
timestamp 1669390400
transform 1 0 49280 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_492
timestamp 1669390400
transform 1 0 56448 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_496
timestamp 1669390400
transform 1 0 56896 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_499
timestamp 1669390400
transform 1 0 57232 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_563
timestamp 1669390400
transform 1 0 64400 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_567
timestamp 1669390400
transform 1 0 64848 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_570
timestamp 1669390400
transform 1 0 65184 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_634
timestamp 1669390400
transform 1 0 72352 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_638
timestamp 1669390400
transform 1 0 72800 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_641
timestamp 1669390400
transform 1 0 73136 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_705
timestamp 1669390400
transform 1 0 80304 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_709
timestamp 1669390400
transform 1 0 80752 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_712
timestamp 1669390400
transform 1 0 81088 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_776
timestamp 1669390400
transform 1 0 88256 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_780
timestamp 1669390400
transform 1 0 88704 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_111_783
timestamp 1669390400
transform 1 0 89040 0 -1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_847
timestamp 1669390400
transform 1 0 96208 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_111_851
timestamp 1669390400
transform 1 0 96656 0 -1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_111_854
timestamp 1669390400
transform 1 0 96992 0 -1 90944
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_111_862
timestamp 1669390400
transform 1 0 97888 0 -1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_112_2
timestamp 1669390400
transform 1 0 1568 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_34
timestamp 1669390400
transform 1 0 5152 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_37
timestamp 1669390400
transform 1 0 5488 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_101
timestamp 1669390400
transform 1 0 12656 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_105
timestamp 1669390400
transform 1 0 13104 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_108
timestamp 1669390400
transform 1 0 13440 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_172
timestamp 1669390400
transform 1 0 20608 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_176
timestamp 1669390400
transform 1 0 21056 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_179
timestamp 1669390400
transform 1 0 21392 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_243
timestamp 1669390400
transform 1 0 28560 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_247
timestamp 1669390400
transform 1 0 29008 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_250
timestamp 1669390400
transform 1 0 29344 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_314
timestamp 1669390400
transform 1 0 36512 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_318
timestamp 1669390400
transform 1 0 36960 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_321
timestamp 1669390400
transform 1 0 37296 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_385
timestamp 1669390400
transform 1 0 44464 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_389
timestamp 1669390400
transform 1 0 44912 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_392
timestamp 1669390400
transform 1 0 45248 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_456
timestamp 1669390400
transform 1 0 52416 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_460
timestamp 1669390400
transform 1 0 52864 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_463
timestamp 1669390400
transform 1 0 53200 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_527
timestamp 1669390400
transform 1 0 60368 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_531
timestamp 1669390400
transform 1 0 60816 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_534
timestamp 1669390400
transform 1 0 61152 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_598
timestamp 1669390400
transform 1 0 68320 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_602
timestamp 1669390400
transform 1 0 68768 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_605
timestamp 1669390400
transform 1 0 69104 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_669
timestamp 1669390400
transform 1 0 76272 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_673
timestamp 1669390400
transform 1 0 76720 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_676
timestamp 1669390400
transform 1 0 77056 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_740
timestamp 1669390400
transform 1 0 84224 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_744
timestamp 1669390400
transform 1 0 84672 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_112_747
timestamp 1669390400
transform 1 0 85008 0 1 90944
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_112_811
timestamp 1669390400
transform 1 0 92176 0 1 90944
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_112_815
timestamp 1669390400
transform 1 0 92624 0 1 90944
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_112_818
timestamp 1669390400
transform 1 0 92960 0 1 90944
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_112_850
timestamp 1669390400
transform 1 0 96544 0 1 90944
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_2
timestamp 1669390400
transform 1 0 1568 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_66
timestamp 1669390400
transform 1 0 8736 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_70
timestamp 1669390400
transform 1 0 9184 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_73
timestamp 1669390400
transform 1 0 9520 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_137
timestamp 1669390400
transform 1 0 16688 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_141
timestamp 1669390400
transform 1 0 17136 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_144
timestamp 1669390400
transform 1 0 17472 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_208
timestamp 1669390400
transform 1 0 24640 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_212
timestamp 1669390400
transform 1 0 25088 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_215
timestamp 1669390400
transform 1 0 25424 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_279
timestamp 1669390400
transform 1 0 32592 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_283
timestamp 1669390400
transform 1 0 33040 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_286
timestamp 1669390400
transform 1 0 33376 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_350
timestamp 1669390400
transform 1 0 40544 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_354
timestamp 1669390400
transform 1 0 40992 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_357
timestamp 1669390400
transform 1 0 41328 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_421
timestamp 1669390400
transform 1 0 48496 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_425
timestamp 1669390400
transform 1 0 48944 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_428
timestamp 1669390400
transform 1 0 49280 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_492
timestamp 1669390400
transform 1 0 56448 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_496
timestamp 1669390400
transform 1 0 56896 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_499
timestamp 1669390400
transform 1 0 57232 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_563
timestamp 1669390400
transform 1 0 64400 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_567
timestamp 1669390400
transform 1 0 64848 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_570
timestamp 1669390400
transform 1 0 65184 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_634
timestamp 1669390400
transform 1 0 72352 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_638
timestamp 1669390400
transform 1 0 72800 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_641
timestamp 1669390400
transform 1 0 73136 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_705
timestamp 1669390400
transform 1 0 80304 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_709
timestamp 1669390400
transform 1 0 80752 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_712
timestamp 1669390400
transform 1 0 81088 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_776
timestamp 1669390400
transform 1 0 88256 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_780
timestamp 1669390400
transform 1 0 88704 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_113_783
timestamp 1669390400
transform 1 0 89040 0 -1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_847
timestamp 1669390400
transform 1 0 96208 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_113_851
timestamp 1669390400
transform 1 0 96656 0 -1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_113_854
timestamp 1669390400
transform 1 0 96992 0 -1 92512
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_113_862
timestamp 1669390400
transform 1 0 97888 0 -1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_114_2
timestamp 1669390400
transform 1 0 1568 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_34
timestamp 1669390400
transform 1 0 5152 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_37
timestamp 1669390400
transform 1 0 5488 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_101
timestamp 1669390400
transform 1 0 12656 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_105
timestamp 1669390400
transform 1 0 13104 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_108
timestamp 1669390400
transform 1 0 13440 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_172
timestamp 1669390400
transform 1 0 20608 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_176
timestamp 1669390400
transform 1 0 21056 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_179
timestamp 1669390400
transform 1 0 21392 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_243
timestamp 1669390400
transform 1 0 28560 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_247
timestamp 1669390400
transform 1 0 29008 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_250
timestamp 1669390400
transform 1 0 29344 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_314
timestamp 1669390400
transform 1 0 36512 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_318
timestamp 1669390400
transform 1 0 36960 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_321
timestamp 1669390400
transform 1 0 37296 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_385
timestamp 1669390400
transform 1 0 44464 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_389
timestamp 1669390400
transform 1 0 44912 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_392
timestamp 1669390400
transform 1 0 45248 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_456
timestamp 1669390400
transform 1 0 52416 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_460
timestamp 1669390400
transform 1 0 52864 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_463
timestamp 1669390400
transform 1 0 53200 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_527
timestamp 1669390400
transform 1 0 60368 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_531
timestamp 1669390400
transform 1 0 60816 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_534
timestamp 1669390400
transform 1 0 61152 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_598
timestamp 1669390400
transform 1 0 68320 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_602
timestamp 1669390400
transform 1 0 68768 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_605
timestamp 1669390400
transform 1 0 69104 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_669
timestamp 1669390400
transform 1 0 76272 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_673
timestamp 1669390400
transform 1 0 76720 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_676
timestamp 1669390400
transform 1 0 77056 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_740
timestamp 1669390400
transform 1 0 84224 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_744
timestamp 1669390400
transform 1 0 84672 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_114_747
timestamp 1669390400
transform 1 0 85008 0 1 92512
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_114_811
timestamp 1669390400
transform 1 0 92176 0 1 92512
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_114_815
timestamp 1669390400
transform 1 0 92624 0 1 92512
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_114_818
timestamp 1669390400
transform 1 0 92960 0 1 92512
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_114_850
timestamp 1669390400
transform 1 0 96544 0 1 92512
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_2
timestamp 1669390400
transform 1 0 1568 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_66
timestamp 1669390400
transform 1 0 8736 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_70
timestamp 1669390400
transform 1 0 9184 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_73
timestamp 1669390400
transform 1 0 9520 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_137
timestamp 1669390400
transform 1 0 16688 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_141
timestamp 1669390400
transform 1 0 17136 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_144
timestamp 1669390400
transform 1 0 17472 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_208
timestamp 1669390400
transform 1 0 24640 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_212
timestamp 1669390400
transform 1 0 25088 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_215
timestamp 1669390400
transform 1 0 25424 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_279
timestamp 1669390400
transform 1 0 32592 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_283
timestamp 1669390400
transform 1 0 33040 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_286
timestamp 1669390400
transform 1 0 33376 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_350
timestamp 1669390400
transform 1 0 40544 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_354
timestamp 1669390400
transform 1 0 40992 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_357
timestamp 1669390400
transform 1 0 41328 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_421
timestamp 1669390400
transform 1 0 48496 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_425
timestamp 1669390400
transform 1 0 48944 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_428
timestamp 1669390400
transform 1 0 49280 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_492
timestamp 1669390400
transform 1 0 56448 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_496
timestamp 1669390400
transform 1 0 56896 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_499
timestamp 1669390400
transform 1 0 57232 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_563
timestamp 1669390400
transform 1 0 64400 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_567
timestamp 1669390400
transform 1 0 64848 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_570
timestamp 1669390400
transform 1 0 65184 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_634
timestamp 1669390400
transform 1 0 72352 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_638
timestamp 1669390400
transform 1 0 72800 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_641
timestamp 1669390400
transform 1 0 73136 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_705
timestamp 1669390400
transform 1 0 80304 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_709
timestamp 1669390400
transform 1 0 80752 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_712
timestamp 1669390400
transform 1 0 81088 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_776
timestamp 1669390400
transform 1 0 88256 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_780
timestamp 1669390400
transform 1 0 88704 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_115_783
timestamp 1669390400
transform 1 0 89040 0 -1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_847
timestamp 1669390400
transform 1 0 96208 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_115_851
timestamp 1669390400
transform 1 0 96656 0 -1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_115_854
timestamp 1669390400
transform 1 0 96992 0 -1 94080
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_115_862
timestamp 1669390400
transform 1 0 97888 0 -1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_2
timestamp 1669390400
transform 1 0 1568 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_34
timestamp 1669390400
transform 1 0 5152 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_37
timestamp 1669390400
transform 1 0 5488 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_101
timestamp 1669390400
transform 1 0 12656 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_105
timestamp 1669390400
transform 1 0 13104 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_108
timestamp 1669390400
transform 1 0 13440 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_172
timestamp 1669390400
transform 1 0 20608 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_176
timestamp 1669390400
transform 1 0 21056 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_179
timestamp 1669390400
transform 1 0 21392 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_243
timestamp 1669390400
transform 1 0 28560 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_247
timestamp 1669390400
transform 1 0 29008 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_250
timestamp 1669390400
transform 1 0 29344 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_314
timestamp 1669390400
transform 1 0 36512 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_318
timestamp 1669390400
transform 1 0 36960 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_321
timestamp 1669390400
transform 1 0 37296 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_385
timestamp 1669390400
transform 1 0 44464 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_389
timestamp 1669390400
transform 1 0 44912 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_392
timestamp 1669390400
transform 1 0 45248 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_456
timestamp 1669390400
transform 1 0 52416 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_460
timestamp 1669390400
transform 1 0 52864 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_463
timestamp 1669390400
transform 1 0 53200 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_527
timestamp 1669390400
transform 1 0 60368 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_531
timestamp 1669390400
transform 1 0 60816 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_534
timestamp 1669390400
transform 1 0 61152 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_598
timestamp 1669390400
transform 1 0 68320 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_602
timestamp 1669390400
transform 1 0 68768 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_605
timestamp 1669390400
transform 1 0 69104 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_669
timestamp 1669390400
transform 1 0 76272 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_673
timestamp 1669390400
transform 1 0 76720 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_676
timestamp 1669390400
transform 1 0 77056 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_740
timestamp 1669390400
transform 1 0 84224 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_744
timestamp 1669390400
transform 1 0 84672 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_116_747
timestamp 1669390400
transform 1 0 85008 0 1 94080
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_116_811
timestamp 1669390400
transform 1 0 92176 0 1 94080
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_116_815
timestamp 1669390400
transform 1 0 92624 0 1 94080
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_116_818
timestamp 1669390400
transform 1 0 92960 0 1 94080
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_116_850
timestamp 1669390400
transform 1 0 96544 0 1 94080
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_2
timestamp 1669390400
transform 1 0 1568 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_66
timestamp 1669390400
transform 1 0 8736 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_70
timestamp 1669390400
transform 1 0 9184 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_73
timestamp 1669390400
transform 1 0 9520 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_137
timestamp 1669390400
transform 1 0 16688 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_141
timestamp 1669390400
transform 1 0 17136 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_144
timestamp 1669390400
transform 1 0 17472 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_208
timestamp 1669390400
transform 1 0 24640 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_212
timestamp 1669390400
transform 1 0 25088 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_215
timestamp 1669390400
transform 1 0 25424 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_279
timestamp 1669390400
transform 1 0 32592 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_283
timestamp 1669390400
transform 1 0 33040 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_286
timestamp 1669390400
transform 1 0 33376 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_350
timestamp 1669390400
transform 1 0 40544 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_354
timestamp 1669390400
transform 1 0 40992 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_357
timestamp 1669390400
transform 1 0 41328 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_421
timestamp 1669390400
transform 1 0 48496 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_425
timestamp 1669390400
transform 1 0 48944 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_428
timestamp 1669390400
transform 1 0 49280 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_492
timestamp 1669390400
transform 1 0 56448 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_496
timestamp 1669390400
transform 1 0 56896 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_499
timestamp 1669390400
transform 1 0 57232 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_563
timestamp 1669390400
transform 1 0 64400 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_567
timestamp 1669390400
transform 1 0 64848 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_570
timestamp 1669390400
transform 1 0 65184 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_634
timestamp 1669390400
transform 1 0 72352 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_638
timestamp 1669390400
transform 1 0 72800 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_641
timestamp 1669390400
transform 1 0 73136 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_705
timestamp 1669390400
transform 1 0 80304 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_709
timestamp 1669390400
transform 1 0 80752 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_712
timestamp 1669390400
transform 1 0 81088 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_776
timestamp 1669390400
transform 1 0 88256 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_780
timestamp 1669390400
transform 1 0 88704 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_117_783
timestamp 1669390400
transform 1 0 89040 0 -1 95648
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_847
timestamp 1669390400
transform 1 0 96208 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_117_851
timestamp 1669390400
transform 1 0 96656 0 -1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_117_854
timestamp 1669390400
transform 1 0 96992 0 -1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_117_862
timestamp 1669390400
transform 1 0 97888 0 -1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_2
timestamp 1669390400
transform 1 0 1568 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_34
timestamp 1669390400
transform 1 0 5152 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_37
timestamp 1669390400
transform 1 0 5488 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_45
timestamp 1669390400
transform 1 0 6384 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_60
timestamp 1669390400
transform 1 0 8064 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_64
timestamp 1669390400
transform 1 0 8512 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_68
timestamp 1669390400
transform 1 0 8960 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_72
timestamp 1669390400
transform 1 0 9408 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_104
timestamp 1669390400
transform 1 0 12992 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_107
timestamp 1669390400
transform 1 0 13328 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_139
timestamp 1669390400
transform 1 0 16912 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_142
timestamp 1669390400
transform 1 0 17248 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_150
timestamp 1669390400
transform 1 0 18144 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_154
timestamp 1669390400
transform 1 0 18592 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_156
timestamp 1669390400
transform 1 0 18816 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_171
timestamp 1669390400
transform 1 0 20496 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_177
timestamp 1669390400
transform 1 0 21168 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_180
timestamp 1669390400
transform 1 0 21504 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_196
timestamp 1669390400
transform 1 0 23296 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_204
timestamp 1669390400
transform 1 0 24192 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_208
timestamp 1669390400
transform 1 0 24640 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_212
timestamp 1669390400
transform 1 0 25088 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_244
timestamp 1669390400
transform 1 0 28672 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_247
timestamp 1669390400
transform 1 0 29008 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_263
timestamp 1669390400
transform 1 0 30800 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_279
timestamp 1669390400
transform 1 0 32592 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_282
timestamp 1669390400
transform 1 0 32928 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_285
timestamp 1669390400
transform 1 0 33264 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_301
timestamp 1669390400
transform 1 0 35056 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_309
timestamp 1669390400
transform 1 0 35952 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_313
timestamp 1669390400
transform 1 0 36400 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_317
timestamp 1669390400
transform 1 0 36848 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_349
timestamp 1669390400
transform 1 0 40432 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_352
timestamp 1669390400
transform 1 0 40768 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_384
timestamp 1669390400
transform 1 0 44352 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_387
timestamp 1669390400
transform 1 0 44688 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_402
timestamp 1669390400
transform 1 0 46368 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_406
timestamp 1669390400
transform 1 0 46816 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_414
timestamp 1669390400
transform 1 0 47712 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_418
timestamp 1669390400
transform 1 0 48160 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_422
timestamp 1669390400
transform 1 0 48608 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_454
timestamp 1669390400
transform 1 0 52192 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_457
timestamp 1669390400
transform 1 0 52528 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_489
timestamp 1669390400
transform 1 0 56112 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_492
timestamp 1669390400
transform 1 0 56448 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_507
timestamp 1669390400
transform 1 0 58128 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_511
timestamp 1669390400
transform 1 0 58576 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_519
timestamp 1669390400
transform 1 0 59472 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_523
timestamp 1669390400
transform 1 0 59920 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_527
timestamp 1669390400
transform 1 0 60368 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_559
timestamp 1669390400
transform 1 0 63952 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_562
timestamp 1669390400
transform 1 0 64288 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_594
timestamp 1669390400
transform 1 0 67872 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_597
timestamp 1669390400
transform 1 0 68208 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_615
timestamp 1669390400
transform 1 0 70224 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_619
timestamp 1669390400
transform 1 0 70672 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_627
timestamp 1669390400
transform 1 0 71568 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_629
timestamp 1669390400
transform 1 0 71792 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_632
timestamp 1669390400
transform 1 0 72128 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_664
timestamp 1669390400
transform 1 0 75712 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_667
timestamp 1669390400
transform 1 0 76048 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_699
timestamp 1669390400
transform 1 0 79632 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_702
timestamp 1669390400
transform 1 0 79968 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_710
timestamp 1669390400
transform 1 0 80864 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_726
timestamp 1669390400
transform 1 0 82656 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_730
timestamp 1669390400
transform 1 0 83104 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_734
timestamp 1669390400
transform 1 0 83552 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_737
timestamp 1669390400
transform 1 0 83888 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_769
timestamp 1669390400
transform 1 0 87472 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_118_772
timestamp 1669390400
transform 1 0 87808 0 1 95648
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_804
timestamp 1669390400
transform 1 0 91392 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_807
timestamp 1669390400
transform 1 0 91728 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_118_815
timestamp 1669390400
transform 1 0 92624 0 1 95648
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_821
timestamp 1669390400
transform 1 0 93296 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_118_837
timestamp 1669390400
transform 1 0 95088 0 1 95648
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_118_839
timestamp 1669390400
transform 1 0 95312 0 1 95648
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_118_842
timestamp 1669390400
transform 1 0 95648 0 1 95648
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_118_858
timestamp 1669390400
transform 1 0 97440 0 1 95648
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 98560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 98560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 98560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 98560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 98560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 98560 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 98560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 98560 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 98560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 98560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 98560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 98560 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 98560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 98560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 98560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 98560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 98560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 98560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 98560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 98560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 98560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 98560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 98560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 98560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 98560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 98560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 98560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 98560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 98560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 98560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 98560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 98560 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 98560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 98560 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 98560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 98560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 98560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 98560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 98560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 98560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 98560 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 98560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 98560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 98560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 98560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 98560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 98560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 98560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 98560 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 98560 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 98560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 98560 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 98560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 98560 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 98560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 98560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 98560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 98560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 98560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 98560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 98560 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 98560 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 98560 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 98560 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 98560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 98560 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 98560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 98560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 98560 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 98560 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 98560 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 98560 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 98560 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1669390400
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1669390400
transform -1 0 98560 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1669390400
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1669390400
transform -1 0 98560 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1669390400
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1669390400
transform -1 0 98560 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1669390400
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1669390400
transform -1 0 98560 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1669390400
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1669390400
transform -1 0 98560 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1669390400
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1669390400
transform -1 0 98560 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1669390400
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1669390400
transform -1 0 98560 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1669390400
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1669390400
transform -1 0 98560 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1669390400
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1669390400
transform -1 0 98560 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1669390400
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1669390400
transform -1 0 98560 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1669390400
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1669390400
transform -1 0 98560 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1669390400
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1669390400
transform -1 0 98560 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1669390400
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1669390400
transform -1 0 98560 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1669390400
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1669390400
transform -1 0 98560 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1669390400
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1669390400
transform -1 0 98560 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1669390400
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1669390400
transform -1 0 98560 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1669390400
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1669390400
transform -1 0 98560 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1669390400
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1669390400
transform -1 0 98560 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1669390400
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1669390400
transform -1 0 98560 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1669390400
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1669390400
transform -1 0 98560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1669390400
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1669390400
transform -1 0 98560 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_188
timestamp 1669390400
transform 1 0 1344 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_189
timestamp 1669390400
transform -1 0 98560 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_190
timestamp 1669390400
transform 1 0 1344 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_191
timestamp 1669390400
transform -1 0 98560 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_192
timestamp 1669390400
transform 1 0 1344 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_193
timestamp 1669390400
transform -1 0 98560 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_194
timestamp 1669390400
transform 1 0 1344 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_195
timestamp 1669390400
transform -1 0 98560 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_196
timestamp 1669390400
transform 1 0 1344 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_197
timestamp 1669390400
transform -1 0 98560 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_198
timestamp 1669390400
transform 1 0 1344 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_199
timestamp 1669390400
transform -1 0 98560 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_200
timestamp 1669390400
transform 1 0 1344 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_201
timestamp 1669390400
transform -1 0 98560 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_202
timestamp 1669390400
transform 1 0 1344 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_203
timestamp 1669390400
transform -1 0 98560 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_204
timestamp 1669390400
transform 1 0 1344 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_205
timestamp 1669390400
transform -1 0 98560 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_206
timestamp 1669390400
transform 1 0 1344 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_207
timestamp 1669390400
transform -1 0 98560 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_208
timestamp 1669390400
transform 1 0 1344 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_209
timestamp 1669390400
transform -1 0 98560 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_210
timestamp 1669390400
transform 1 0 1344 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_211
timestamp 1669390400
transform -1 0 98560 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_212
timestamp 1669390400
transform 1 0 1344 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_213
timestamp 1669390400
transform -1 0 98560 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_214
timestamp 1669390400
transform 1 0 1344 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_215
timestamp 1669390400
transform -1 0 98560 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_216
timestamp 1669390400
transform 1 0 1344 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_217
timestamp 1669390400
transform -1 0 98560 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_218
timestamp 1669390400
transform 1 0 1344 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_219
timestamp 1669390400
transform -1 0 98560 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_220
timestamp 1669390400
transform 1 0 1344 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_221
timestamp 1669390400
transform -1 0 98560 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_222
timestamp 1669390400
transform 1 0 1344 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_223
timestamp 1669390400
transform -1 0 98560 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_224
timestamp 1669390400
transform 1 0 1344 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_225
timestamp 1669390400
transform -1 0 98560 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_226
timestamp 1669390400
transform 1 0 1344 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_227
timestamp 1669390400
transform -1 0 98560 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_228
timestamp 1669390400
transform 1 0 1344 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_229
timestamp 1669390400
transform -1 0 98560 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_230
timestamp 1669390400
transform 1 0 1344 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_231
timestamp 1669390400
transform -1 0 98560 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_232
timestamp 1669390400
transform 1 0 1344 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_233
timestamp 1669390400
transform -1 0 98560 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_234
timestamp 1669390400
transform 1 0 1344 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_235
timestamp 1669390400
transform -1 0 98560 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_236
timestamp 1669390400
transform 1 0 1344 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_237
timestamp 1669390400
transform -1 0 98560 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 84784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 92736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 80864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 88816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 96768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 84784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 92736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 80864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 88816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 96768 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 84784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 92736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 80864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 88816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 96768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 84784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 92736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 80864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 88816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 96768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 84784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 92736 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 80864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 88816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 96768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 84784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 92736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 80864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 88816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 96768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1669390400
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1669390400
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1669390400
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1669390400
transform 1 0 84784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1669390400
transform 1 0 92736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1669390400
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1669390400
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1669390400
transform 1 0 80864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1669390400
transform 1 0 88816 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1669390400
transform 1 0 96768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1669390400
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1669390400
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1669390400
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1669390400
transform 1 0 84784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1669390400
transform 1 0 92736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1669390400
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1669390400
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1669390400
transform 1 0 80864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1669390400
transform 1 0 88816 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1669390400
transform 1 0 96768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1669390400
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1669390400
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1669390400
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1669390400
transform 1 0 84784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1669390400
transform 1 0 92736 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1669390400
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1669390400
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1669390400
transform 1 0 80864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1669390400
transform 1 0 88816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1669390400
transform 1 0 96768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1669390400
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1669390400
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1669390400
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1669390400
transform 1 0 84784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1669390400
transform 1 0 92736 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1669390400
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1669390400
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1669390400
transform 1 0 80864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1669390400
transform 1 0 88816 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1669390400
transform 1 0 96768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1669390400
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1669390400
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1669390400
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1669390400
transform 1 0 84784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1669390400
transform 1 0 92736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1669390400
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1669390400
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1669390400
transform 1 0 80864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1669390400
transform 1 0 88816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1669390400
transform 1 0 96768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1669390400
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1669390400
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1669390400
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1669390400
transform 1 0 84784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1669390400
transform 1 0 92736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1669390400
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1669390400
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1669390400
transform 1 0 80864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1669390400
transform 1 0 88816 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1669390400
transform 1 0 96768 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1669390400
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1669390400
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1669390400
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1669390400
transform 1 0 84784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1669390400
transform 1 0 92736 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1669390400
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1669390400
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1669390400
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1669390400
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1669390400
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1669390400
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1669390400
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1669390400
transform 1 0 80864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1669390400
transform 1 0 88816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1669390400
transform 1 0 96768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1669390400
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1669390400
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1669390400
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1669390400
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1669390400
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1669390400
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1669390400
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1669390400
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1669390400
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1669390400
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1669390400
transform 1 0 84784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1669390400
transform 1 0 92736 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1669390400
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1669390400
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1669390400
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1669390400
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1669390400
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1669390400
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1669390400
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1669390400
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1669390400
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1669390400
transform 1 0 80864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1669390400
transform 1 0 88816 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1669390400
transform 1 0 96768 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1669390400
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1669390400
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1669390400
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1669390400
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1669390400
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1669390400
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1669390400
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1669390400
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1669390400
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1669390400
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1100
timestamp 1669390400
transform 1 0 84784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1101
timestamp 1669390400
transform 1 0 92736 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1102
timestamp 1669390400
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1103
timestamp 1669390400
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1104
timestamp 1669390400
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1105
timestamp 1669390400
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1106
timestamp 1669390400
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1107
timestamp 1669390400
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1108
timestamp 1669390400
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1109
timestamp 1669390400
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1110
timestamp 1669390400
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1111
timestamp 1669390400
transform 1 0 80864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1112
timestamp 1669390400
transform 1 0 88816 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1113
timestamp 1669390400
transform 1 0 96768 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1114
timestamp 1669390400
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1115
timestamp 1669390400
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1116
timestamp 1669390400
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1117
timestamp 1669390400
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1118
timestamp 1669390400
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1119
timestamp 1669390400
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1120
timestamp 1669390400
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1121
timestamp 1669390400
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1122
timestamp 1669390400
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1123
timestamp 1669390400
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1124
timestamp 1669390400
transform 1 0 84784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1125
timestamp 1669390400
transform 1 0 92736 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1126
timestamp 1669390400
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1127
timestamp 1669390400
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1128
timestamp 1669390400
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1129
timestamp 1669390400
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1130
timestamp 1669390400
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1131
timestamp 1669390400
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1132
timestamp 1669390400
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1133
timestamp 1669390400
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1134
timestamp 1669390400
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1135
timestamp 1669390400
transform 1 0 80864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1136
timestamp 1669390400
transform 1 0 88816 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1137
timestamp 1669390400
transform 1 0 96768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1138
timestamp 1669390400
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1139
timestamp 1669390400
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1140
timestamp 1669390400
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1141
timestamp 1669390400
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1142
timestamp 1669390400
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1143
timestamp 1669390400
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1144
timestamp 1669390400
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1145
timestamp 1669390400
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1146
timestamp 1669390400
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1147
timestamp 1669390400
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1148
timestamp 1669390400
transform 1 0 84784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1149
timestamp 1669390400
transform 1 0 92736 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1150
timestamp 1669390400
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1151
timestamp 1669390400
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1152
timestamp 1669390400
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1153
timestamp 1669390400
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1154
timestamp 1669390400
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1155
timestamp 1669390400
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1156
timestamp 1669390400
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1157
timestamp 1669390400
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1158
timestamp 1669390400
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1159
timestamp 1669390400
transform 1 0 80864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1160
timestamp 1669390400
transform 1 0 88816 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1161
timestamp 1669390400
transform 1 0 96768 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1162
timestamp 1669390400
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1163
timestamp 1669390400
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1164
timestamp 1669390400
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1165
timestamp 1669390400
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1166
timestamp 1669390400
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1167
timestamp 1669390400
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1168
timestamp 1669390400
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1169
timestamp 1669390400
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1170
timestamp 1669390400
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1171
timestamp 1669390400
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1172
timestamp 1669390400
transform 1 0 84784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1173
timestamp 1669390400
transform 1 0 92736 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1174
timestamp 1669390400
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1175
timestamp 1669390400
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1176
timestamp 1669390400
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1177
timestamp 1669390400
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1178
timestamp 1669390400
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1179
timestamp 1669390400
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1180
timestamp 1669390400
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1181
timestamp 1669390400
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1182
timestamp 1669390400
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1183
timestamp 1669390400
transform 1 0 80864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1184
timestamp 1669390400
transform 1 0 88816 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1185
timestamp 1669390400
transform 1 0 96768 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1186
timestamp 1669390400
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1187
timestamp 1669390400
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1188
timestamp 1669390400
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1189
timestamp 1669390400
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1190
timestamp 1669390400
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1191
timestamp 1669390400
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1192
timestamp 1669390400
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1193
timestamp 1669390400
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1194
timestamp 1669390400
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1195
timestamp 1669390400
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1196
timestamp 1669390400
transform 1 0 84784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1197
timestamp 1669390400
transform 1 0 92736 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1198
timestamp 1669390400
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1199
timestamp 1669390400
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1200
timestamp 1669390400
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1201
timestamp 1669390400
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1202
timestamp 1669390400
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1203
timestamp 1669390400
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1204
timestamp 1669390400
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1205
timestamp 1669390400
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1206
timestamp 1669390400
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1207
timestamp 1669390400
transform 1 0 80864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1208
timestamp 1669390400
transform 1 0 88816 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1209
timestamp 1669390400
transform 1 0 96768 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1210
timestamp 1669390400
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1211
timestamp 1669390400
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1212
timestamp 1669390400
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1213
timestamp 1669390400
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1214
timestamp 1669390400
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1215
timestamp 1669390400
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1216
timestamp 1669390400
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1217
timestamp 1669390400
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1218
timestamp 1669390400
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1219
timestamp 1669390400
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1220
timestamp 1669390400
transform 1 0 84784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1221
timestamp 1669390400
transform 1 0 92736 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1222
timestamp 1669390400
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1223
timestamp 1669390400
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1224
timestamp 1669390400
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1225
timestamp 1669390400
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1226
timestamp 1669390400
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1227
timestamp 1669390400
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1228
timestamp 1669390400
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1229
timestamp 1669390400
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1230
timestamp 1669390400
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1231
timestamp 1669390400
transform 1 0 80864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1232
timestamp 1669390400
transform 1 0 88816 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1233
timestamp 1669390400
transform 1 0 96768 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1234
timestamp 1669390400
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1235
timestamp 1669390400
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1236
timestamp 1669390400
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1237
timestamp 1669390400
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1238
timestamp 1669390400
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1239
timestamp 1669390400
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1240
timestamp 1669390400
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1241
timestamp 1669390400
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1242
timestamp 1669390400
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1243
timestamp 1669390400
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1244
timestamp 1669390400
transform 1 0 84784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1245
timestamp 1669390400
transform 1 0 92736 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1246
timestamp 1669390400
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1247
timestamp 1669390400
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1248
timestamp 1669390400
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1249
timestamp 1669390400
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1250
timestamp 1669390400
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1251
timestamp 1669390400
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1252
timestamp 1669390400
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1253
timestamp 1669390400
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1254
timestamp 1669390400
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1255
timestamp 1669390400
transform 1 0 80864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1256
timestamp 1669390400
transform 1 0 88816 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1257
timestamp 1669390400
transform 1 0 96768 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1258
timestamp 1669390400
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1259
timestamp 1669390400
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1260
timestamp 1669390400
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1261
timestamp 1669390400
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1262
timestamp 1669390400
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1263
timestamp 1669390400
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1264
timestamp 1669390400
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1265
timestamp 1669390400
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1266
timestamp 1669390400
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1267
timestamp 1669390400
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1268
timestamp 1669390400
transform 1 0 84784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1269
timestamp 1669390400
transform 1 0 92736 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1270
timestamp 1669390400
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1271
timestamp 1669390400
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1272
timestamp 1669390400
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1273
timestamp 1669390400
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1274
timestamp 1669390400
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1275
timestamp 1669390400
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1276
timestamp 1669390400
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1277
timestamp 1669390400
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1278
timestamp 1669390400
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1279
timestamp 1669390400
transform 1 0 80864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1280
timestamp 1669390400
transform 1 0 88816 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1281
timestamp 1669390400
transform 1 0 96768 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1282
timestamp 1669390400
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1283
timestamp 1669390400
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1284
timestamp 1669390400
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1285
timestamp 1669390400
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1286
timestamp 1669390400
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1287
timestamp 1669390400
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1288
timestamp 1669390400
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1289
timestamp 1669390400
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1290
timestamp 1669390400
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1291
timestamp 1669390400
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1292
timestamp 1669390400
transform 1 0 84784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1293
timestamp 1669390400
transform 1 0 92736 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1294
timestamp 1669390400
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1295
timestamp 1669390400
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1296
timestamp 1669390400
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1297
timestamp 1669390400
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1298
timestamp 1669390400
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1299
timestamp 1669390400
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1300
timestamp 1669390400
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1301
timestamp 1669390400
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1302
timestamp 1669390400
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1303
timestamp 1669390400
transform 1 0 80864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1304
timestamp 1669390400
transform 1 0 88816 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1305
timestamp 1669390400
transform 1 0 96768 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1306
timestamp 1669390400
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1307
timestamp 1669390400
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1308
timestamp 1669390400
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1309
timestamp 1669390400
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1310
timestamp 1669390400
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1311
timestamp 1669390400
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1312
timestamp 1669390400
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1313
timestamp 1669390400
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1314
timestamp 1669390400
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1315
timestamp 1669390400
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1316
timestamp 1669390400
transform 1 0 84784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1317
timestamp 1669390400
transform 1 0 92736 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1318
timestamp 1669390400
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1319
timestamp 1669390400
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1320
timestamp 1669390400
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1321
timestamp 1669390400
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1322
timestamp 1669390400
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1323
timestamp 1669390400
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1324
timestamp 1669390400
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1325
timestamp 1669390400
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1326
timestamp 1669390400
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1327
timestamp 1669390400
transform 1 0 80864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1328
timestamp 1669390400
transform 1 0 88816 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1329
timestamp 1669390400
transform 1 0 96768 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1330
timestamp 1669390400
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1331
timestamp 1669390400
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1332
timestamp 1669390400
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1333
timestamp 1669390400
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1334
timestamp 1669390400
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1335
timestamp 1669390400
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1336
timestamp 1669390400
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1337
timestamp 1669390400
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1338
timestamp 1669390400
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1339
timestamp 1669390400
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1340
timestamp 1669390400
transform 1 0 84784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1341
timestamp 1669390400
transform 1 0 92736 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1342
timestamp 1669390400
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1343
timestamp 1669390400
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1344
timestamp 1669390400
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1345
timestamp 1669390400
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1346
timestamp 1669390400
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1347
timestamp 1669390400
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1348
timestamp 1669390400
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1349
timestamp 1669390400
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1350
timestamp 1669390400
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1351
timestamp 1669390400
transform 1 0 80864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1352
timestamp 1669390400
transform 1 0 88816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1353
timestamp 1669390400
transform 1 0 96768 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1354
timestamp 1669390400
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1355
timestamp 1669390400
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1356
timestamp 1669390400
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1357
timestamp 1669390400
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1358
timestamp 1669390400
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1359
timestamp 1669390400
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1360
timestamp 1669390400
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1361
timestamp 1669390400
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1362
timestamp 1669390400
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1363
timestamp 1669390400
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1364
timestamp 1669390400
transform 1 0 84784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1365
timestamp 1669390400
transform 1 0 92736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1366
timestamp 1669390400
transform 1 0 9296 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1367
timestamp 1669390400
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1368
timestamp 1669390400
transform 1 0 25200 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1369
timestamp 1669390400
transform 1 0 33152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1370
timestamp 1669390400
transform 1 0 41104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1371
timestamp 1669390400
transform 1 0 49056 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1372
timestamp 1669390400
transform 1 0 57008 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1373
timestamp 1669390400
transform 1 0 64960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1374
timestamp 1669390400
transform 1 0 72912 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1375
timestamp 1669390400
transform 1 0 80864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1376
timestamp 1669390400
transform 1 0 88816 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1377
timestamp 1669390400
transform 1 0 96768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1378
timestamp 1669390400
transform 1 0 5264 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1379
timestamp 1669390400
transform 1 0 13216 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1380
timestamp 1669390400
transform 1 0 21168 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1381
timestamp 1669390400
transform 1 0 29120 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1382
timestamp 1669390400
transform 1 0 37072 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1383
timestamp 1669390400
transform 1 0 45024 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1384
timestamp 1669390400
transform 1 0 52976 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1385
timestamp 1669390400
transform 1 0 60928 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1386
timestamp 1669390400
transform 1 0 68880 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1387
timestamp 1669390400
transform 1 0 76832 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1388
timestamp 1669390400
transform 1 0 84784 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1389
timestamp 1669390400
transform 1 0 92736 0 1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1390
timestamp 1669390400
transform 1 0 9296 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1391
timestamp 1669390400
transform 1 0 17248 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1392
timestamp 1669390400
transform 1 0 25200 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1393
timestamp 1669390400
transform 1 0 33152 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1394
timestamp 1669390400
transform 1 0 41104 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1395
timestamp 1669390400
transform 1 0 49056 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1396
timestamp 1669390400
transform 1 0 57008 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1397
timestamp 1669390400
transform 1 0 64960 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1398
timestamp 1669390400
transform 1 0 72912 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1399
timestamp 1669390400
transform 1 0 80864 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1400
timestamp 1669390400
transform 1 0 88816 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1401
timestamp 1669390400
transform 1 0 96768 0 -1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1402
timestamp 1669390400
transform 1 0 5264 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1403
timestamp 1669390400
transform 1 0 13216 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1404
timestamp 1669390400
transform 1 0 21168 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1405
timestamp 1669390400
transform 1 0 29120 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1406
timestamp 1669390400
transform 1 0 37072 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1407
timestamp 1669390400
transform 1 0 45024 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1408
timestamp 1669390400
transform 1 0 52976 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1409
timestamp 1669390400
transform 1 0 60928 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1410
timestamp 1669390400
transform 1 0 68880 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1411
timestamp 1669390400
transform 1 0 76832 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1412
timestamp 1669390400
transform 1 0 84784 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1413
timestamp 1669390400
transform 1 0 92736 0 1 78400
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1414
timestamp 1669390400
transform 1 0 9296 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1415
timestamp 1669390400
transform 1 0 17248 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1416
timestamp 1669390400
transform 1 0 25200 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1417
timestamp 1669390400
transform 1 0 33152 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1418
timestamp 1669390400
transform 1 0 41104 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1419
timestamp 1669390400
transform 1 0 49056 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1420
timestamp 1669390400
transform 1 0 57008 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1421
timestamp 1669390400
transform 1 0 64960 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1422
timestamp 1669390400
transform 1 0 72912 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1423
timestamp 1669390400
transform 1 0 80864 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1424
timestamp 1669390400
transform 1 0 88816 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1425
timestamp 1669390400
transform 1 0 96768 0 -1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1426
timestamp 1669390400
transform 1 0 5264 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1427
timestamp 1669390400
transform 1 0 13216 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1428
timestamp 1669390400
transform 1 0 21168 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1429
timestamp 1669390400
transform 1 0 29120 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1430
timestamp 1669390400
transform 1 0 37072 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1431
timestamp 1669390400
transform 1 0 45024 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1432
timestamp 1669390400
transform 1 0 52976 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1433
timestamp 1669390400
transform 1 0 60928 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1434
timestamp 1669390400
transform 1 0 68880 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1435
timestamp 1669390400
transform 1 0 76832 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1436
timestamp 1669390400
transform 1 0 84784 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1437
timestamp 1669390400
transform 1 0 92736 0 1 79968
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1438
timestamp 1669390400
transform 1 0 9296 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1439
timestamp 1669390400
transform 1 0 17248 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1440
timestamp 1669390400
transform 1 0 25200 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1441
timestamp 1669390400
transform 1 0 33152 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1442
timestamp 1669390400
transform 1 0 41104 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1443
timestamp 1669390400
transform 1 0 49056 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1444
timestamp 1669390400
transform 1 0 57008 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1445
timestamp 1669390400
transform 1 0 64960 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1446
timestamp 1669390400
transform 1 0 72912 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1447
timestamp 1669390400
transform 1 0 80864 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1448
timestamp 1669390400
transform 1 0 88816 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1449
timestamp 1669390400
transform 1 0 96768 0 -1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1450
timestamp 1669390400
transform 1 0 5264 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1451
timestamp 1669390400
transform 1 0 13216 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1452
timestamp 1669390400
transform 1 0 21168 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1453
timestamp 1669390400
transform 1 0 29120 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1454
timestamp 1669390400
transform 1 0 37072 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1455
timestamp 1669390400
transform 1 0 45024 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1456
timestamp 1669390400
transform 1 0 52976 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1457
timestamp 1669390400
transform 1 0 60928 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1458
timestamp 1669390400
transform 1 0 68880 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1459
timestamp 1669390400
transform 1 0 76832 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1460
timestamp 1669390400
transform 1 0 84784 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1461
timestamp 1669390400
transform 1 0 92736 0 1 81536
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1462
timestamp 1669390400
transform 1 0 9296 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1463
timestamp 1669390400
transform 1 0 17248 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1464
timestamp 1669390400
transform 1 0 25200 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1465
timestamp 1669390400
transform 1 0 33152 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1466
timestamp 1669390400
transform 1 0 41104 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1467
timestamp 1669390400
transform 1 0 49056 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1468
timestamp 1669390400
transform 1 0 57008 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1469
timestamp 1669390400
transform 1 0 64960 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1470
timestamp 1669390400
transform 1 0 72912 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1471
timestamp 1669390400
transform 1 0 80864 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1472
timestamp 1669390400
transform 1 0 88816 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1473
timestamp 1669390400
transform 1 0 96768 0 -1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1474
timestamp 1669390400
transform 1 0 5264 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1475
timestamp 1669390400
transform 1 0 13216 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1476
timestamp 1669390400
transform 1 0 21168 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1477
timestamp 1669390400
transform 1 0 29120 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1478
timestamp 1669390400
transform 1 0 37072 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1479
timestamp 1669390400
transform 1 0 45024 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1480
timestamp 1669390400
transform 1 0 52976 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1481
timestamp 1669390400
transform 1 0 60928 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1482
timestamp 1669390400
transform 1 0 68880 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1483
timestamp 1669390400
transform 1 0 76832 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1484
timestamp 1669390400
transform 1 0 84784 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1485
timestamp 1669390400
transform 1 0 92736 0 1 83104
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1486
timestamp 1669390400
transform 1 0 9296 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1487
timestamp 1669390400
transform 1 0 17248 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1488
timestamp 1669390400
transform 1 0 25200 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1489
timestamp 1669390400
transform 1 0 33152 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1490
timestamp 1669390400
transform 1 0 41104 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1491
timestamp 1669390400
transform 1 0 49056 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1492
timestamp 1669390400
transform 1 0 57008 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1493
timestamp 1669390400
transform 1 0 64960 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1494
timestamp 1669390400
transform 1 0 72912 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1495
timestamp 1669390400
transform 1 0 80864 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1496
timestamp 1669390400
transform 1 0 88816 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1497
timestamp 1669390400
transform 1 0 96768 0 -1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1498
timestamp 1669390400
transform 1 0 5264 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1499
timestamp 1669390400
transform 1 0 13216 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1500
timestamp 1669390400
transform 1 0 21168 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1501
timestamp 1669390400
transform 1 0 29120 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1502
timestamp 1669390400
transform 1 0 37072 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1503
timestamp 1669390400
transform 1 0 45024 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1504
timestamp 1669390400
transform 1 0 52976 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1505
timestamp 1669390400
transform 1 0 60928 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1506
timestamp 1669390400
transform 1 0 68880 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1507
timestamp 1669390400
transform 1 0 76832 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1508
timestamp 1669390400
transform 1 0 84784 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1509
timestamp 1669390400
transform 1 0 92736 0 1 84672
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1510
timestamp 1669390400
transform 1 0 9296 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1511
timestamp 1669390400
transform 1 0 17248 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1512
timestamp 1669390400
transform 1 0 25200 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1513
timestamp 1669390400
transform 1 0 33152 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1514
timestamp 1669390400
transform 1 0 41104 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1515
timestamp 1669390400
transform 1 0 49056 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1516
timestamp 1669390400
transform 1 0 57008 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1517
timestamp 1669390400
transform 1 0 64960 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1518
timestamp 1669390400
transform 1 0 72912 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1519
timestamp 1669390400
transform 1 0 80864 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1520
timestamp 1669390400
transform 1 0 88816 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1521
timestamp 1669390400
transform 1 0 96768 0 -1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1522
timestamp 1669390400
transform 1 0 5264 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1523
timestamp 1669390400
transform 1 0 13216 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1524
timestamp 1669390400
transform 1 0 21168 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1525
timestamp 1669390400
transform 1 0 29120 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1526
timestamp 1669390400
transform 1 0 37072 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1527
timestamp 1669390400
transform 1 0 45024 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1528
timestamp 1669390400
transform 1 0 52976 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1529
timestamp 1669390400
transform 1 0 60928 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1530
timestamp 1669390400
transform 1 0 68880 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1531
timestamp 1669390400
transform 1 0 76832 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1532
timestamp 1669390400
transform 1 0 84784 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1533
timestamp 1669390400
transform 1 0 92736 0 1 86240
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1534
timestamp 1669390400
transform 1 0 9296 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1535
timestamp 1669390400
transform 1 0 17248 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1536
timestamp 1669390400
transform 1 0 25200 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1537
timestamp 1669390400
transform 1 0 33152 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1538
timestamp 1669390400
transform 1 0 41104 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1539
timestamp 1669390400
transform 1 0 49056 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1540
timestamp 1669390400
transform 1 0 57008 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1541
timestamp 1669390400
transform 1 0 64960 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1542
timestamp 1669390400
transform 1 0 72912 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1543
timestamp 1669390400
transform 1 0 80864 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1544
timestamp 1669390400
transform 1 0 88816 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1545
timestamp 1669390400
transform 1 0 96768 0 -1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1546
timestamp 1669390400
transform 1 0 5264 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1547
timestamp 1669390400
transform 1 0 13216 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1548
timestamp 1669390400
transform 1 0 21168 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1549
timestamp 1669390400
transform 1 0 29120 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1550
timestamp 1669390400
transform 1 0 37072 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1551
timestamp 1669390400
transform 1 0 45024 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1552
timestamp 1669390400
transform 1 0 52976 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1553
timestamp 1669390400
transform 1 0 60928 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1554
timestamp 1669390400
transform 1 0 68880 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1555
timestamp 1669390400
transform 1 0 76832 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1556
timestamp 1669390400
transform 1 0 84784 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1557
timestamp 1669390400
transform 1 0 92736 0 1 87808
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1558
timestamp 1669390400
transform 1 0 9296 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1559
timestamp 1669390400
transform 1 0 17248 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1560
timestamp 1669390400
transform 1 0 25200 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1561
timestamp 1669390400
transform 1 0 33152 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1562
timestamp 1669390400
transform 1 0 41104 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1563
timestamp 1669390400
transform 1 0 49056 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1564
timestamp 1669390400
transform 1 0 57008 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1565
timestamp 1669390400
transform 1 0 64960 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1566
timestamp 1669390400
transform 1 0 72912 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1567
timestamp 1669390400
transform 1 0 80864 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1568
timestamp 1669390400
transform 1 0 88816 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1569
timestamp 1669390400
transform 1 0 96768 0 -1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1570
timestamp 1669390400
transform 1 0 5264 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1571
timestamp 1669390400
transform 1 0 13216 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1572
timestamp 1669390400
transform 1 0 21168 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1573
timestamp 1669390400
transform 1 0 29120 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1574
timestamp 1669390400
transform 1 0 37072 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1575
timestamp 1669390400
transform 1 0 45024 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1576
timestamp 1669390400
transform 1 0 52976 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1577
timestamp 1669390400
transform 1 0 60928 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1578
timestamp 1669390400
transform 1 0 68880 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1579
timestamp 1669390400
transform 1 0 76832 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1580
timestamp 1669390400
transform 1 0 84784 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1581
timestamp 1669390400
transform 1 0 92736 0 1 89376
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1582
timestamp 1669390400
transform 1 0 9296 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1583
timestamp 1669390400
transform 1 0 17248 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1584
timestamp 1669390400
transform 1 0 25200 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1585
timestamp 1669390400
transform 1 0 33152 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1586
timestamp 1669390400
transform 1 0 41104 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1587
timestamp 1669390400
transform 1 0 49056 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1588
timestamp 1669390400
transform 1 0 57008 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1589
timestamp 1669390400
transform 1 0 64960 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1590
timestamp 1669390400
transform 1 0 72912 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1591
timestamp 1669390400
transform 1 0 80864 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1592
timestamp 1669390400
transform 1 0 88816 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1593
timestamp 1669390400
transform 1 0 96768 0 -1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1594
timestamp 1669390400
transform 1 0 5264 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1595
timestamp 1669390400
transform 1 0 13216 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1596
timestamp 1669390400
transform 1 0 21168 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1597
timestamp 1669390400
transform 1 0 29120 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1598
timestamp 1669390400
transform 1 0 37072 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1599
timestamp 1669390400
transform 1 0 45024 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1600
timestamp 1669390400
transform 1 0 52976 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1601
timestamp 1669390400
transform 1 0 60928 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1602
timestamp 1669390400
transform 1 0 68880 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1603
timestamp 1669390400
transform 1 0 76832 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1604
timestamp 1669390400
transform 1 0 84784 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1605
timestamp 1669390400
transform 1 0 92736 0 1 90944
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1606
timestamp 1669390400
transform 1 0 9296 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1607
timestamp 1669390400
transform 1 0 17248 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1608
timestamp 1669390400
transform 1 0 25200 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1609
timestamp 1669390400
transform 1 0 33152 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1610
timestamp 1669390400
transform 1 0 41104 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1611
timestamp 1669390400
transform 1 0 49056 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1612
timestamp 1669390400
transform 1 0 57008 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1613
timestamp 1669390400
transform 1 0 64960 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1614
timestamp 1669390400
transform 1 0 72912 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1615
timestamp 1669390400
transform 1 0 80864 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1616
timestamp 1669390400
transform 1 0 88816 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1617
timestamp 1669390400
transform 1 0 96768 0 -1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1618
timestamp 1669390400
transform 1 0 5264 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1619
timestamp 1669390400
transform 1 0 13216 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1620
timestamp 1669390400
transform 1 0 21168 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1621
timestamp 1669390400
transform 1 0 29120 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1622
timestamp 1669390400
transform 1 0 37072 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1623
timestamp 1669390400
transform 1 0 45024 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1624
timestamp 1669390400
transform 1 0 52976 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1625
timestamp 1669390400
transform 1 0 60928 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1626
timestamp 1669390400
transform 1 0 68880 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1627
timestamp 1669390400
transform 1 0 76832 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1628
timestamp 1669390400
transform 1 0 84784 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1629
timestamp 1669390400
transform 1 0 92736 0 1 92512
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1630
timestamp 1669390400
transform 1 0 9296 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1631
timestamp 1669390400
transform 1 0 17248 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1632
timestamp 1669390400
transform 1 0 25200 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1633
timestamp 1669390400
transform 1 0 33152 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1634
timestamp 1669390400
transform 1 0 41104 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1635
timestamp 1669390400
transform 1 0 49056 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1636
timestamp 1669390400
transform 1 0 57008 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1637
timestamp 1669390400
transform 1 0 64960 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1638
timestamp 1669390400
transform 1 0 72912 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1639
timestamp 1669390400
transform 1 0 80864 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1640
timestamp 1669390400
transform 1 0 88816 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1641
timestamp 1669390400
transform 1 0 96768 0 -1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1642
timestamp 1669390400
transform 1 0 5264 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1643
timestamp 1669390400
transform 1 0 13216 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1644
timestamp 1669390400
transform 1 0 21168 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1645
timestamp 1669390400
transform 1 0 29120 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1646
timestamp 1669390400
transform 1 0 37072 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1647
timestamp 1669390400
transform 1 0 45024 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1648
timestamp 1669390400
transform 1 0 52976 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1649
timestamp 1669390400
transform 1 0 60928 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1650
timestamp 1669390400
transform 1 0 68880 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1651
timestamp 1669390400
transform 1 0 76832 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1652
timestamp 1669390400
transform 1 0 84784 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1653
timestamp 1669390400
transform 1 0 92736 0 1 94080
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1654
timestamp 1669390400
transform 1 0 9296 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1655
timestamp 1669390400
transform 1 0 17248 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1656
timestamp 1669390400
transform 1 0 25200 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1657
timestamp 1669390400
transform 1 0 33152 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1658
timestamp 1669390400
transform 1 0 41104 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1659
timestamp 1669390400
transform 1 0 49056 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1660
timestamp 1669390400
transform 1 0 57008 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1661
timestamp 1669390400
transform 1 0 64960 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1662
timestamp 1669390400
transform 1 0 72912 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1663
timestamp 1669390400
transform 1 0 80864 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1664
timestamp 1669390400
transform 1 0 88816 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1665
timestamp 1669390400
transform 1 0 96768 0 -1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1666
timestamp 1669390400
transform 1 0 5264 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1667
timestamp 1669390400
transform 1 0 9184 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1668
timestamp 1669390400
transform 1 0 13104 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1669
timestamp 1669390400
transform 1 0 17024 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1670
timestamp 1669390400
transform 1 0 20944 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1671
timestamp 1669390400
transform 1 0 24864 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1672
timestamp 1669390400
transform 1 0 28784 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1673
timestamp 1669390400
transform 1 0 32704 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1674
timestamp 1669390400
transform 1 0 36624 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1675
timestamp 1669390400
transform 1 0 40544 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1676
timestamp 1669390400
transform 1 0 44464 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1677
timestamp 1669390400
transform 1 0 48384 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1678
timestamp 1669390400
transform 1 0 52304 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1679
timestamp 1669390400
transform 1 0 56224 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1680
timestamp 1669390400
transform 1 0 60144 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1681
timestamp 1669390400
transform 1 0 64064 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1682
timestamp 1669390400
transform 1 0 67984 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1683
timestamp 1669390400
transform 1 0 71904 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1684
timestamp 1669390400
transform 1 0 75824 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1685
timestamp 1669390400
transform 1 0 79744 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1686
timestamp 1669390400
transform 1 0 83664 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1687
timestamp 1669390400
transform 1 0 87584 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1688
timestamp 1669390400
transform 1 0 91504 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1689
timestamp 1669390400
transform 1 0 95424 0 1 95648
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0831_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 71904 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0832_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 77952 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0833_
timestamp 1669390400
transform 1 0 78624 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0834_
timestamp 1669390400
transform 1 0 78064 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0835_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 78848 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0836_
timestamp 1669390400
transform 1 0 68096 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0837_
timestamp 1669390400
transform 1 0 69328 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0838_
timestamp 1669390400
transform 1 0 78736 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0839_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 77168 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0840_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 80640 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0841_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 72576 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0842_
timestamp 1669390400
transform -1 0 79856 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0843_
timestamp 1669390400
transform -1 0 82992 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0844_
timestamp 1669390400
transform -1 0 76608 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0845_
timestamp 1669390400
transform 1 0 66416 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0846_
timestamp 1669390400
transform 1 0 78288 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0847_
timestamp 1669390400
transform 1 0 79184 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0848_
timestamp 1669390400
transform 1 0 69664 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0849_
timestamp 1669390400
transform 1 0 70448 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0850_
timestamp 1669390400
transform 1 0 79744 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0851_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 81200 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0852_
timestamp 1669390400
transform -1 0 80416 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0853_
timestamp 1669390400
transform 1 0 73248 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0854_
timestamp 1669390400
transform 1 0 75600 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0855_
timestamp 1669390400
transform -1 0 72128 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0856_
timestamp 1669390400
transform 1 0 75376 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0857_
timestamp 1669390400
transform 1 0 77168 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0858_
timestamp 1669390400
transform 1 0 79408 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0859_
timestamp 1669390400
transform 1 0 78848 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0860_
timestamp 1669390400
transform 1 0 70336 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0861_
timestamp 1669390400
transform 1 0 71456 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0862_
timestamp 1669390400
transform 1 0 80080 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0863_
timestamp 1669390400
transform 1 0 79296 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0864_
timestamp 1669390400
transform 1 0 70896 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0865_
timestamp 1669390400
transform 1 0 70000 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0866_
timestamp 1669390400
transform 1 0 79296 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0867_
timestamp 1669390400
transform 1 0 80192 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0868_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 81424 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0869_
timestamp 1669390400
transform 1 0 85120 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0870_
timestamp 1669390400
transform -1 0 85680 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0871_
timestamp 1669390400
transform 1 0 89152 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0872_
timestamp 1669390400
transform -1 0 86800 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0873_
timestamp 1669390400
transform -1 0 88816 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0874_
timestamp 1669390400
transform -1 0 84448 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0875_
timestamp 1669390400
transform 1 0 84672 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0876_
timestamp 1669390400
transform -1 0 84336 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0877_
timestamp 1669390400
transform 1 0 85680 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0878_
timestamp 1669390400
transform -1 0 78288 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0879_
timestamp 1669390400
transform -1 0 72352 0 -1 78400
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0880_
timestamp 1669390400
transform 1 0 85120 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0881_
timestamp 1669390400
transform -1 0 84448 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0882_
timestamp 1669390400
transform 1 0 78288 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0883_
timestamp 1669390400
transform 1 0 89152 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0884_
timestamp 1669390400
transform -1 0 86800 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0885_
timestamp 1669390400
transform 1 0 85904 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0886_
timestamp 1669390400
transform -1 0 85344 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0887_
timestamp 1669390400
transform -1 0 81984 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0888_
timestamp 1669390400
transform -1 0 72128 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0889_
timestamp 1669390400
transform 1 0 83552 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0890_
timestamp 1669390400
transform -1 0 84112 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0891_
timestamp 1669390400
transform 1 0 85904 0 -1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0892_
timestamp 1669390400
transform 1 0 85120 0 -1 81536
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0893_
timestamp 1669390400
transform -1 0 87024 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0894_
timestamp 1669390400
transform 1 0 87920 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0895_
timestamp 1669390400
transform -1 0 88032 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0896_
timestamp 1669390400
transform 1 0 81200 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0897_
timestamp 1669390400
transform -1 0 84896 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0898_
timestamp 1669390400
transform -1 0 78400 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0899_
timestamp 1669390400
transform 1 0 85120 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0900_
timestamp 1669390400
transform -1 0 86016 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0901_
timestamp 1669390400
transform -1 0 83664 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1669390400
transform -1 0 68208 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0903_
timestamp 1669390400
transform 1 0 66304 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0904_
timestamp 1669390400
transform 1 0 69216 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0905_
timestamp 1669390400
transform -1 0 69888 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0906_
timestamp 1669390400
transform 1 0 66976 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0907_
timestamp 1669390400
transform 1 0 66528 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0908_
timestamp 1669390400
transform -1 0 71008 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0909_
timestamp 1669390400
transform 1 0 67872 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0910_
timestamp 1669390400
transform -1 0 72464 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0911_
timestamp 1669390400
transform -1 0 71344 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0912_
timestamp 1669390400
transform 1 0 69664 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0913_
timestamp 1669390400
transform -1 0 71792 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0914_
timestamp 1669390400
transform -1 0 67760 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0915_
timestamp 1669390400
transform -1 0 69104 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0916_
timestamp 1669390400
transform -1 0 70336 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0917_
timestamp 1669390400
transform -1 0 68208 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0918_
timestamp 1669390400
transform 1 0 67312 0 1 65856
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0919_
timestamp 1669390400
transform 1 0 57344 0 -1 79968
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0920_
timestamp 1669390400
transform 1 0 58464 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0921_
timestamp 1669390400
transform 1 0 57344 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0922_
timestamp 1669390400
transform -1 0 58240 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0923_
timestamp 1669390400
transform -1 0 61376 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0924_
timestamp 1669390400
transform 1 0 59024 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0925_
timestamp 1669390400
transform -1 0 66080 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0926_
timestamp 1669390400
transform -1 0 63728 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0927_
timestamp 1669390400
transform -1 0 60256 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0928_
timestamp 1669390400
transform 1 0 57232 0 1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0929_
timestamp 1669390400
transform -1 0 60816 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0930_
timestamp 1669390400
transform 1 0 77168 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0931_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 72800 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0932_
timestamp 1669390400
transform 1 0 53312 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0933_
timestamp 1669390400
transform 1 0 57344 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0934_
timestamp 1669390400
transform -1 0 58576 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0935_
timestamp 1669390400
transform -1 0 59472 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0936_
timestamp 1669390400
transform 1 0 61712 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0937_
timestamp 1669390400
transform 1 0 61712 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0938_
timestamp 1669390400
transform -1 0 57120 0 1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0939_
timestamp 1669390400
transform 1 0 59136 0 -1 78400
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0940_
timestamp 1669390400
transform -1 0 59136 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0941_
timestamp 1669390400
transform 1 0 53536 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0942_
timestamp 1669390400
transform 1 0 57344 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0943_
timestamp 1669390400
transform 1 0 54432 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0944_
timestamp 1669390400
transform 1 0 54880 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _0945_
timestamp 1669390400
transform 1 0 61264 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0946_
timestamp 1669390400
transform 1 0 61824 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0947_
timestamp 1669390400
transform -1 0 59024 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0948_
timestamp 1669390400
transform 1 0 81984 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0949_
timestamp 1669390400
transform -1 0 71680 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0950_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 72352 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0951_
timestamp 1669390400
transform 1 0 74816 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0952_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 76160 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0953_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 74592 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0954_
timestamp 1669390400
transform -1 0 73808 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0955_
timestamp 1669390400
transform 1 0 77616 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0956_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 81984 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0957_
timestamp 1669390400
transform 1 0 81088 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0958_
timestamp 1669390400
transform 1 0 77168 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0959_
timestamp 1669390400
transform -1 0 79296 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0960_
timestamp 1669390400
transform 1 0 83104 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0961_
timestamp 1669390400
transform -1 0 84448 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0962_
timestamp 1669390400
transform -1 0 84672 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0963_
timestamp 1669390400
transform 1 0 85120 0 1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0964_
timestamp 1669390400
transform 1 0 85120 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0965_
timestamp 1669390400
transform 1 0 81648 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0966_
timestamp 1669390400
transform 1 0 67872 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0967_
timestamp 1669390400
transform 1 0 81760 0 1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0968_
timestamp 1669390400
transform 1 0 81312 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0969_
timestamp 1669390400
transform -1 0 84672 0 1 56448
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0970_
timestamp 1669390400
transform 1 0 85120 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0971_
timestamp 1669390400
transform 1 0 66192 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0972_
timestamp 1669390400
transform 1 0 65968 0 -1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0973_
timestamp 1669390400
transform -1 0 65856 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0974_
timestamp 1669390400
transform 1 0 85120 0 1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0975_
timestamp 1669390400
transform 1 0 82768 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0976_
timestamp 1669390400
transform 1 0 48272 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0977_
timestamp 1669390400
transform -1 0 67760 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0978_
timestamp 1669390400
transform 1 0 49168 0 1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0979_
timestamp 1669390400
transform 1 0 48272 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0980_
timestamp 1669390400
transform 1 0 65408 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0981_
timestamp 1669390400
transform 1 0 64176 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0982_
timestamp 1669390400
transform 1 0 48272 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0983_
timestamp 1669390400
transform 1 0 49168 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0984_
timestamp 1669390400
transform 1 0 48272 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0985_
timestamp 1669390400
transform 1 0 49504 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0986_
timestamp 1669390400
transform 1 0 47376 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0987_
timestamp 1669390400
transform -1 0 52304 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0988_
timestamp 1669390400
transform 1 0 74816 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0989_
timestamp 1669390400
transform 1 0 49392 0 -1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0990_
timestamp 1669390400
transform 1 0 48272 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0991_
timestamp 1669390400
transform 1 0 51520 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0992_
timestamp 1669390400
transform 1 0 47712 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0993_
timestamp 1669390400
transform 1 0 49616 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0994_
timestamp 1669390400
transform 1 0 49168 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0995_
timestamp 1669390400
transform 1 0 93744 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0996_
timestamp 1669390400
transform 1 0 70784 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0997_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 75040 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0998_
timestamp 1669390400
transform 1 0 75040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _0999_
timestamp 1669390400
transform -1 0 96656 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1000_
timestamp 1669390400
transform -1 0 97776 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1001_
timestamp 1669390400
transform 1 0 77168 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1002_
timestamp 1669390400
transform 1 0 76608 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1003_
timestamp 1669390400
transform 1 0 90048 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1004_
timestamp 1669390400
transform 1 0 89152 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1005_
timestamp 1669390400
transform -1 0 89824 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1006_
timestamp 1669390400
transform -1 0 96656 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1007_
timestamp 1669390400
transform 1 0 95648 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1008_
timestamp 1669390400
transform 1 0 82880 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1009_
timestamp 1669390400
transform 1 0 71568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1010_
timestamp 1669390400
transform 1 0 82656 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1011_
timestamp 1669390400
transform -1 0 82432 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1012_
timestamp 1669390400
transform 1 0 85568 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1013_
timestamp 1669390400
transform -1 0 86128 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1014_
timestamp 1669390400
transform 1 0 69216 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1015_
timestamp 1669390400
transform 1 0 69440 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1016_
timestamp 1669390400
transform -1 0 68768 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1017_
timestamp 1669390400
transform 1 0 82992 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1018_
timestamp 1669390400
transform 1 0 82096 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1019_
timestamp 1669390400
transform 1 0 57344 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1020_
timestamp 1669390400
transform -1 0 70112 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1021_
timestamp 1669390400
transform 1 0 61936 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1022_
timestamp 1669390400
transform -1 0 60144 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1023_
timestamp 1669390400
transform 1 0 69664 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1024_
timestamp 1669390400
transform -1 0 67872 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1025_
timestamp 1669390400
transform 1 0 54208 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1026_
timestamp 1669390400
transform 1 0 58352 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1027_
timestamp 1669390400
transform 1 0 57456 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1028_
timestamp 1669390400
transform 1 0 63168 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1029_
timestamp 1669390400
transform -1 0 60368 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1030_
timestamp 1669390400
transform 1 0 50960 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1031_
timestamp 1669390400
transform -1 0 71120 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1032_
timestamp 1669390400
transform 1 0 49504 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1033_
timestamp 1669390400
transform 1 0 48272 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1034_
timestamp 1669390400
transform 1 0 57344 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1035_
timestamp 1669390400
transform -1 0 56784 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1036_
timestamp 1669390400
transform -1 0 75264 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1037_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 69888 0 1 61152
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1038_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 71568 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1039_
timestamp 1669390400
transform 1 0 72464 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1040_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 73024 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1041_
timestamp 1669390400
transform 1 0 74928 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1042_
timestamp 1669390400
transform 1 0 74144 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1043_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 74144 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1044_
timestamp 1669390400
transform 1 0 74144 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1045_
timestamp 1669390400
transform 1 0 75824 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1046_
timestamp 1669390400
transform -1 0 75152 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1047_
timestamp 1669390400
transform 1 0 51408 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1048_
timestamp 1669390400
transform -1 0 51408 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1049_
timestamp 1669390400
transform 1 0 81200 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1050_
timestamp 1669390400
transform -1 0 75488 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1051_
timestamp 1669390400
transform 1 0 77168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1052_
timestamp 1669390400
transform 1 0 94976 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1053_
timestamp 1669390400
transform 1 0 93632 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1054_
timestamp 1669390400
transform 1 0 78736 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1055_
timestamp 1669390400
transform 1 0 78848 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1056_
timestamp 1669390400
transform -1 0 92288 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1057_
timestamp 1669390400
transform -1 0 93296 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1058_
timestamp 1669390400
transform -1 0 96656 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1059_
timestamp 1669390400
transform -1 0 97776 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1060_
timestamp 1669390400
transform -1 0 75712 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1061_
timestamp 1669390400
transform 1 0 87024 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1062_
timestamp 1669390400
transform -1 0 84112 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1063_
timestamp 1669390400
transform 1 0 89152 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1064_
timestamp 1669390400
transform 1 0 88928 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1065_
timestamp 1669390400
transform 1 0 73248 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1066_
timestamp 1669390400
transform -1 0 71344 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1067_
timestamp 1669390400
transform 1 0 85344 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1068_
timestamp 1669390400
transform 1 0 84000 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1069_
timestamp 1669390400
transform -1 0 74256 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1070_
timestamp 1669390400
transform 1 0 61488 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1071_
timestamp 1669390400
transform 1 0 60144 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1072_
timestamp 1669390400
transform 1 0 71568 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1073_
timestamp 1669390400
transform -1 0 72240 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1074_
timestamp 1669390400
transform -1 0 63392 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1075_
timestamp 1669390400
transform 1 0 60144 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1076_
timestamp 1669390400
transform 1 0 64736 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1077_
timestamp 1669390400
transform -1 0 65968 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1078_
timestamp 1669390400
transform 1 0 75264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1079_
timestamp 1669390400
transform -1 0 64848 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1080_
timestamp 1669390400
transform -1 0 65968 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1081_
timestamp 1669390400
transform 1 0 63168 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1082_
timestamp 1669390400
transform -1 0 64512 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1083_
timestamp 1669390400
transform 1 0 70672 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1084_
timestamp 1669390400
transform 1 0 69776 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1085_
timestamp 1669390400
transform 1 0 63168 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1086_
timestamp 1669390400
transform 1 0 62272 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1087_
timestamp 1669390400
transform 1 0 93072 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1088_
timestamp 1669390400
transform 1 0 71904 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1089_
timestamp 1669390400
transform -1 0 73024 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1090_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 76720 0 1 54880
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1091_
timestamp 1669390400
transform 1 0 77168 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1092_
timestamp 1669390400
transform 1 0 95312 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1093_
timestamp 1669390400
transform 1 0 70112 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1094_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 73248 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1095_
timestamp 1669390400
transform 1 0 75712 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1096_
timestamp 1669390400
transform 1 0 95984 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1097_
timestamp 1669390400
transform -1 0 97664 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1098_
timestamp 1669390400
transform -1 0 81760 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1099_
timestamp 1669390400
transform 1 0 78960 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1100_
timestamp 1669390400
transform 1 0 79744 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1101_
timestamp 1669390400
transform 1 0 90944 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1102_
timestamp 1669390400
transform -1 0 95088 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1103_
timestamp 1669390400
transform -1 0 97664 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1104_
timestamp 1669390400
transform 1 0 92960 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1105_
timestamp 1669390400
transform 1 0 74592 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1106_
timestamp 1669390400
transform 1 0 93856 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1107_
timestamp 1669390400
transform 1 0 95200 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1108_
timestamp 1669390400
transform 1 0 89712 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1109_
timestamp 1669390400
transform 1 0 93856 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1110_
timestamp 1669390400
transform 1 0 95984 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1111_
timestamp 1669390400
transform -1 0 96656 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1112_
timestamp 1669390400
transform 1 0 93072 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1113_
timestamp 1669390400
transform -1 0 93632 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1114_
timestamp 1669390400
transform 1 0 67872 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1115_
timestamp 1669390400
transform -1 0 73920 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1116_
timestamp 1669390400
transform 1 0 68208 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1117_
timestamp 1669390400
transform -1 0 74816 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1118_
timestamp 1669390400
transform -1 0 72576 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1119_
timestamp 1669390400
transform -1 0 70224 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1120_
timestamp 1669390400
transform 1 0 94416 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1121_
timestamp 1669390400
transform -1 0 97664 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1122_
timestamp 1669390400
transform 1 0 56224 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1123_
timestamp 1669390400
transform 1 0 62384 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1124_
timestamp 1669390400
transform -1 0 66752 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1125_
timestamp 1669390400
transform -1 0 65856 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1126_
timestamp 1669390400
transform -1 0 73808 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1127_
timestamp 1669390400
transform -1 0 72464 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1128_
timestamp 1669390400
transform 1 0 55104 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1129_
timestamp 1669390400
transform -1 0 62160 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1130_
timestamp 1669390400
transform -1 0 65856 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1131_
timestamp 1669390400
transform 1 0 60480 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1132_
timestamp 1669390400
transform 1 0 74704 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1133_
timestamp 1669390400
transform -1 0 66640 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1669390400
transform -1 0 65296 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1135_
timestamp 1669390400
transform 1 0 51408 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1136_
timestamp 1669390400
transform 1 0 61264 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1137_
timestamp 1669390400
transform -1 0 66640 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1138_
timestamp 1669390400
transform -1 0 64512 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1139_
timestamp 1669390400
transform -1 0 64288 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1140_
timestamp 1669390400
transform -1 0 63728 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1141_
timestamp 1669390400
transform 1 0 75936 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1142_
timestamp 1669390400
transform 1 0 75040 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1143_
timestamp 1669390400
transform 1 0 74368 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1144_
timestamp 1669390400
transform 1 0 65184 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1145_
timestamp 1669390400
transform -1 0 65856 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1146_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 77168 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1147_
timestamp 1669390400
transform 1 0 77952 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1148_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 75264 0 -1 58016
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1149_
timestamp 1669390400
transform 1 0 79856 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1150_
timestamp 1669390400
transform 1 0 94192 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1151_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 76272 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1152_
timestamp 1669390400
transform 1 0 78400 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1153_
timestamp 1669390400
transform 1 0 97104 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1154_
timestamp 1669390400
transform -1 0 95088 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1155_
timestamp 1669390400
transform -1 0 82096 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1156_
timestamp 1669390400
transform 1 0 80192 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1157_
timestamp 1669390400
transform 1 0 81200 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1158_
timestamp 1669390400
transform 1 0 92624 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1159_
timestamp 1669390400
transform -1 0 96656 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1160_
timestamp 1669390400
transform 1 0 92624 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1161_
timestamp 1669390400
transform -1 0 79520 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1162_
timestamp 1669390400
transform 1 0 96880 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1163_
timestamp 1669390400
transform -1 0 98224 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1164_
timestamp 1669390400
transform 1 0 93408 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1165_
timestamp 1669390400
transform -1 0 96096 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1166_
timestamp 1669390400
transform -1 0 95872 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1167_
timestamp 1669390400
transform -1 0 94528 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1168_
timestamp 1669390400
transform 1 0 92064 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1169_
timestamp 1669390400
transform -1 0 75040 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1170_
timestamp 1669390400
transform -1 0 67984 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1171_
timestamp 1669390400
transform -1 0 69888 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1172_
timestamp 1669390400
transform -1 0 68544 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1173_
timestamp 1669390400
transform -1 0 67760 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1174_
timestamp 1669390400
transform -1 0 95312 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1175_
timestamp 1669390400
transform -1 0 94752 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1176_
timestamp 1669390400
transform 1 0 56224 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1177_
timestamp 1669390400
transform -1 0 57904 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1178_
timestamp 1669390400
transform -1 0 57904 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1179_
timestamp 1669390400
transform -1 0 69552 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1180_
timestamp 1669390400
transform -1 0 68208 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1181_
timestamp 1669390400
transform 1 0 56224 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1182_
timestamp 1669390400
transform -1 0 58464 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1183_
timestamp 1669390400
transform -1 0 57904 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1184_
timestamp 1669390400
transform 1 0 77168 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1185_
timestamp 1669390400
transform -1 0 58688 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1186_
timestamp 1669390400
transform 1 0 54208 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1187_
timestamp 1669390400
transform -1 0 56000 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1188_
timestamp 1669390400
transform -1 0 57680 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1189_
timestamp 1669390400
transform 1 0 52864 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1190_
timestamp 1669390400
transform -1 0 57568 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1191_
timestamp 1669390400
transform -1 0 55776 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1192_
timestamp 1669390400
transform 1 0 77168 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1193_
timestamp 1669390400
transform 1 0 76608 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1194_
timestamp 1669390400
transform 1 0 78064 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1195_
timestamp 1669390400
transform 1 0 56000 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1196_
timestamp 1669390400
transform -1 0 58688 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1197_
timestamp 1669390400
transform -1 0 94304 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1198_
timestamp 1669390400
transform 1 0 75488 0 -1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1199_
timestamp 1669390400
transform 1 0 73584 0 -1 62720
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1200_
timestamp 1669390400
transform 1 0 75824 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1201_
timestamp 1669390400
transform 1 0 96544 0 1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1202_
timestamp 1669390400
transform -1 0 96096 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1203_
timestamp 1669390400
transform -1 0 79632 0 -1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1204_
timestamp 1669390400
transform -1 0 78736 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1205_
timestamp 1669390400
transform 1 0 93072 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1206_
timestamp 1669390400
transform 1 0 93184 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1207_
timestamp 1669390400
transform 1 0 93072 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1208_
timestamp 1669390400
transform 1 0 94976 0 -1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1209_
timestamp 1669390400
transform -1 0 97776 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1210_
timestamp 1669390400
transform -1 0 89824 0 -1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1211_
timestamp 1669390400
transform -1 0 74144 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1212_
timestamp 1669390400
transform 1 0 89152 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1213_
timestamp 1669390400
transform 1 0 88032 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1214_
timestamp 1669390400
transform 1 0 91168 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1215_
timestamp 1669390400
transform -1 0 90832 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1216_
timestamp 1669390400
transform 1 0 68096 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1217_
timestamp 1669390400
transform 1 0 70336 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1218_
timestamp 1669390400
transform -1 0 69888 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1219_
timestamp 1669390400
transform 1 0 89152 0 -1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1220_
timestamp 1669390400
transform -1 0 88704 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1221_
timestamp 1669390400
transform 1 0 53424 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1222_
timestamp 1669390400
transform -1 0 72464 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1223_
timestamp 1669390400
transform 1 0 57792 0 1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1224_
timestamp 1669390400
transform -1 0 56560 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1225_
timestamp 1669390400
transform 1 0 69216 0 1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1226_
timestamp 1669390400
transform -1 0 68768 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1227_
timestamp 1669390400
transform -1 0 55664 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1228_
timestamp 1669390400
transform 1 0 55888 0 1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1229_
timestamp 1669390400
transform -1 0 55664 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1230_
timestamp 1669390400
transform 1 0 58352 0 1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1231_
timestamp 1669390400
transform 1 0 56000 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1232_
timestamp 1669390400
transform -1 0 51968 0 -1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1233_
timestamp 1669390400
transform 1 0 73696 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1234_
timestamp 1669390400
transform 1 0 49952 0 -1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1235_
timestamp 1669390400
transform 1 0 47712 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1236_
timestamp 1669390400
transform 1 0 57344 0 -1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1237_
timestamp 1669390400
transform -1 0 54768 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1238_
timestamp 1669390400
transform 1 0 78064 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1239_
timestamp 1669390400
transform 1 0 79296 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1240_
timestamp 1669390400
transform 1 0 50176 0 -1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1241_
timestamp 1669390400
transform 1 0 49504 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1242_
timestamp 1669390400
transform -1 0 77728 0 -1 59584
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1243_
timestamp 1669390400
transform 1 0 77168 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1244_
timestamp 1669390400
transform -1 0 96656 0 -1 78400
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1245_
timestamp 1669390400
transform -1 0 97776 0 -1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1246_
timestamp 1669390400
transform -1 0 79520 0 -1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1247_
timestamp 1669390400
transform 1 0 77616 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1248_
timestamp 1669390400
transform 1 0 94976 0 -1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1249_
timestamp 1669390400
transform 1 0 95424 0 -1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1250_
timestamp 1669390400
transform 1 0 94976 0 -1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1251_
timestamp 1669390400
transform -1 0 96320 0 -1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1252_
timestamp 1669390400
transform 1 0 73248 0 -1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1253_
timestamp 1669390400
transform 1 0 90944 0 1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1254_
timestamp 1669390400
transform 1 0 91392 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1255_
timestamp 1669390400
transform 1 0 94976 0 1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1256_
timestamp 1669390400
transform 1 0 95424 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1257_
timestamp 1669390400
transform 1 0 71120 0 -1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1258_
timestamp 1669390400
transform -1 0 70784 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1259_
timestamp 1669390400
transform 1 0 90944 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1260_
timestamp 1669390400
transform -1 0 93744 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1261_
timestamp 1669390400
transform -1 0 73920 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1262_
timestamp 1669390400
transform 1 0 57792 0 -1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1263_
timestamp 1669390400
transform -1 0 57904 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1264_
timestamp 1669390400
transform 1 0 71120 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1265_
timestamp 1669390400
transform -1 0 68768 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1266_
timestamp 1669390400
transform 1 0 61264 0 1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1267_
timestamp 1669390400
transform -1 0 61936 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1268_
timestamp 1669390400
transform -1 0 60032 0 1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1269_
timestamp 1669390400
transform -1 0 60368 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1270_
timestamp 1669390400
transform 1 0 74144 0 1 86240
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1271_
timestamp 1669390400
transform 1 0 65968 0 1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1272_
timestamp 1669390400
transform -1 0 63952 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1273_
timestamp 1669390400
transform 1 0 63168 0 -1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1274_
timestamp 1669390400
transform 1 0 61264 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1275_
timestamp 1669390400
transform -1 0 75376 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1276_
timestamp 1669390400
transform 1 0 74592 0 1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1277_
timestamp 1669390400
transform 1 0 74592 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1278_
timestamp 1669390400
transform 1 0 63168 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1279_
timestamp 1669390400
transform 1 0 63392 0 1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1280_
timestamp 1669390400
transform 1 0 73584 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1281_
timestamp 1669390400
transform 1 0 74704 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1282_
timestamp 1669390400
transform 1 0 92624 0 -1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1283_
timestamp 1669390400
transform 1 0 93072 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1284_
timestamp 1669390400
transform -1 0 78848 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1285_
timestamp 1669390400
transform -1 0 76608 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1286_
timestamp 1669390400
transform 1 0 93072 0 1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1287_
timestamp 1669390400
transform 1 0 93072 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1288_
timestamp 1669390400
transform 1 0 93744 0 -1 79968
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1289_
timestamp 1669390400
transform 1 0 91392 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1290_
timestamp 1669390400
transform 1 0 72464 0 1 83104
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1291_
timestamp 1669390400
transform 1 0 87360 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1292_
timestamp 1669390400
transform 1 0 86800 0 -1 87808
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1293_
timestamp 1669390400
transform 1 0 88032 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1294_
timestamp 1669390400
transform -1 0 89824 0 -1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1295_
timestamp 1669390400
transform 1 0 69888 0 -1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1296_
timestamp 1669390400
transform -1 0 69888 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1297_
timestamp 1669390400
transform 1 0 88592 0 1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1298_
timestamp 1669390400
transform -1 0 86688 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1299_
timestamp 1669390400
transform -1 0 72688 0 -1 84672
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1300_
timestamp 1669390400
transform 1 0 52976 0 -1 87808
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1301_
timestamp 1669390400
transform -1 0 52752 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1302_
timestamp 1669390400
transform 1 0 69216 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1303_
timestamp 1669390400
transform -1 0 68544 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1304_
timestamp 1669390400
transform 1 0 55216 0 -1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1305_
timestamp 1669390400
transform -1 0 55888 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1306_
timestamp 1669390400
transform 1 0 53312 0 1 86240
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1307_
timestamp 1669390400
transform -1 0 52752 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1308_
timestamp 1669390400
transform 1 0 72688 0 1 81536
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1309_
timestamp 1669390400
transform -1 0 63952 0 -1 79968
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1310_
timestamp 1669390400
transform -1 0 64512 0 -1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1311_
timestamp 1669390400
transform 1 0 58352 0 1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1312_
timestamp 1669390400
transform 1 0 57680 0 1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1313_
timestamp 1669390400
transform 1 0 74704 0 1 84672
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1314_
timestamp 1669390400
transform -1 0 75936 0 1 86240
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1315_
timestamp 1669390400
transform 1 0 62048 0 1 81536
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1316_
timestamp 1669390400
transform -1 0 62160 0 -1 83104
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1317_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 71456 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1318_
timestamp 1669390400
transform 1 0 72240 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1319_
timestamp 1669390400
transform 1 0 75152 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1320_
timestamp 1669390400
transform 1 0 96544 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1321_
timestamp 1669390400
transform -1 0 92624 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1322_
timestamp 1669390400
transform 1 0 74592 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1323_
timestamp 1669390400
transform -1 0 77840 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1324_
timestamp 1669390400
transform 1 0 90048 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1325_
timestamp 1669390400
transform 1 0 89152 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1326_
timestamp 1669390400
transform -1 0 92624 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1327_
timestamp 1669390400
transform 1 0 93072 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1328_
timestamp 1669390400
transform 1 0 71120 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1329_
timestamp 1669390400
transform 1 0 81536 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1330_
timestamp 1669390400
transform -1 0 81872 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1331_
timestamp 1669390400
transform 1 0 81872 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1332_
timestamp 1669390400
transform 1 0 81536 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1333_
timestamp 1669390400
transform 1 0 69216 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1334_
timestamp 1669390400
transform -1 0 68544 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1335_
timestamp 1669390400
transform 1 0 82096 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1336_
timestamp 1669390400
transform -1 0 80080 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1337_
timestamp 1669390400
transform -1 0 70448 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1338_
timestamp 1669390400
transform -1 0 59360 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1339_
timestamp 1669390400
transform 1 0 59360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1340_
timestamp 1669390400
transform 1 0 66976 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1341_
timestamp 1669390400
transform -1 0 66752 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1342_
timestamp 1669390400
transform 1 0 56112 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1343_
timestamp 1669390400
transform -1 0 56000 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1344_
timestamp 1669390400
transform 1 0 57456 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1345_
timestamp 1669390400
transform 1 0 56224 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1346_
timestamp 1669390400
transform 1 0 71568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1347_
timestamp 1669390400
transform 1 0 51184 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1348_
timestamp 1669390400
transform 1 0 49392 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1349_
timestamp 1669390400
transform 1 0 55216 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1350_
timestamp 1669390400
transform -1 0 55552 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1351_
timestamp 1669390400
transform 1 0 74032 0 1 83104
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1352_
timestamp 1669390400
transform 1 0 73808 0 1 84672
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1353_
timestamp 1669390400
transform 1 0 52864 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1354_
timestamp 1669390400
transform -1 0 50960 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1355_
timestamp 1669390400
transform -1 0 78064 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1356_
timestamp 1669390400
transform 1 0 70896 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1357_
timestamp 1669390400
transform 1 0 73248 0 -1 64288
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1358_
timestamp 1669390400
transform 1 0 75040 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1359_
timestamp 1669390400
transform -1 0 94528 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1360_
timestamp 1669390400
transform -1 0 78064 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1361_
timestamp 1669390400
transform -1 0 71344 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1362_
timestamp 1669390400
transform 1 0 75040 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1363_
timestamp 1669390400
transform 1 0 75936 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1364_
timestamp 1669390400
transform -1 0 91056 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1365_
timestamp 1669390400
transform 1 0 89600 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1366_
timestamp 1669390400
transform -1 0 78624 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1367_
timestamp 1669390400
transform 1 0 75376 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1368_
timestamp 1669390400
transform 1 0 76160 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1369_
timestamp 1669390400
transform -1 0 92064 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1370_
timestamp 1669390400
transform -1 0 91280 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1371_
timestamp 1669390400
transform -1 0 90496 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1372_
timestamp 1669390400
transform 1 0 70112 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1373_
timestamp 1669390400
transform 1 0 87360 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1374_
timestamp 1669390400
transform 1 0 88144 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1375_
timestamp 1669390400
transform -1 0 90272 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1376_
timestamp 1669390400
transform -1 0 93184 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1377_
timestamp 1669390400
transform 1 0 89152 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1378_
timestamp 1669390400
transform 1 0 85456 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1379_
timestamp 1669390400
transform 1 0 86240 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1380_
timestamp 1669390400
transform -1 0 69888 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1381_
timestamp 1669390400
transform 1 0 67760 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1382_
timestamp 1669390400
transform -1 0 75936 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1383_
timestamp 1669390400
transform -1 0 70560 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1384_
timestamp 1669390400
transform -1 0 68768 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1385_
timestamp 1669390400
transform -1 0 84112 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1386_
timestamp 1669390400
transform -1 0 83328 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1387_
timestamp 1669390400
transform -1 0 57904 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1388_
timestamp 1669390400
transform -1 0 59472 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1389_
timestamp 1669390400
transform -1 0 56784 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1390_
timestamp 1669390400
transform -1 0 69776 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1391_
timestamp 1669390400
transform -1 0 68656 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1392_
timestamp 1669390400
transform -1 0 55440 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1393_
timestamp 1669390400
transform -1 0 53872 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1394_
timestamp 1669390400
transform -1 0 53872 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1395_
timestamp 1669390400
transform 1 0 71008 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1396_
timestamp 1669390400
transform 1 0 57344 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1397_
timestamp 1669390400
transform 1 0 58128 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1398_
timestamp 1669390400
transform -1 0 53872 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1399_
timestamp 1669390400
transform -1 0 54432 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1400_
timestamp 1669390400
transform -1 0 53648 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1401_
timestamp 1669390400
transform 1 0 54096 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1402_
timestamp 1669390400
transform -1 0 55216 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1403_
timestamp 1669390400
transform 1 0 73248 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1404_
timestamp 1669390400
transform -1 0 73920 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1405_
timestamp 1669390400
transform -1 0 54656 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1406_
timestamp 1669390400
transform -1 0 52864 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1407_
timestamp 1669390400
transform 1 0 72576 0 1 62720
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1408_
timestamp 1669390400
transform 1 0 76272 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1409_
timestamp 1669390400
transform 1 0 88032 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1410_
timestamp 1669390400
transform 1 0 71344 0 1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1411_
timestamp 1669390400
transform 1 0 76160 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1412_
timestamp 1669390400
transform -1 0 90832 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1413_
timestamp 1669390400
transform 1 0 88144 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1414_
timestamp 1669390400
transform -1 0 79296 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1415_
timestamp 1669390400
transform 1 0 78176 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1416_
timestamp 1669390400
transform 1 0 78624 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1417_
timestamp 1669390400
transform -1 0 90608 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1418_
timestamp 1669390400
transform -1 0 89824 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1419_
timestamp 1669390400
transform 1 0 89152 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1420_
timestamp 1669390400
transform 1 0 70448 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1421_
timestamp 1669390400
transform 1 0 87584 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1422_
timestamp 1669390400
transform 1 0 88144 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1423_
timestamp 1669390400
transform -1 0 91392 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1424_
timestamp 1669390400
transform -1 0 93632 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1669390400
transform 1 0 89488 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1426_
timestamp 1669390400
transform 1 0 86800 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1427_
timestamp 1669390400
transform 1 0 87248 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1428_
timestamp 1669390400
transform -1 0 69664 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1429_
timestamp 1669390400
transform 1 0 67648 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1430_
timestamp 1669390400
transform -1 0 72352 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1431_
timestamp 1669390400
transform -1 0 69776 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1432_
timestamp 1669390400
transform -1 0 68768 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1433_
timestamp 1669390400
transform 1 0 88368 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1434_
timestamp 1669390400
transform 1 0 89376 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1435_
timestamp 1669390400
transform 1 0 62384 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1436_
timestamp 1669390400
transform -1 0 65856 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1437_
timestamp 1669390400
transform -1 0 64512 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1438_
timestamp 1669390400
transform -1 0 70560 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1439_
timestamp 1669390400
transform 1 0 66864 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1440_
timestamp 1669390400
transform -1 0 60256 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1441_
timestamp 1669390400
transform -1 0 65856 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1442_
timestamp 1669390400
transform -1 0 62608 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1443_
timestamp 1669390400
transform -1 0 75936 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1444_
timestamp 1669390400
transform -1 0 65296 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1445_
timestamp 1669390400
transform -1 0 63392 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1446_
timestamp 1669390400
transform -1 0 62160 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1447_
timestamp 1669390400
transform -1 0 63728 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1448_
timestamp 1669390400
transform 1 0 60704 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1449_
timestamp 1669390400
transform -1 0 66080 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1450_
timestamp 1669390400
transform -1 0 60816 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1451_
timestamp 1669390400
transform -1 0 76608 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1452_
timestamp 1669390400
transform -1 0 76160 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1453_
timestamp 1669390400
transform -1 0 65856 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1454_
timestamp 1669390400
transform -1 0 64176 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1455_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 74816 0 1 61152
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1456_
timestamp 1669390400
transform 1 0 75600 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1457_
timestamp 1669390400
transform 1 0 94976 0 -1 64288
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1669390400
transform 1 0 94080 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1459_
timestamp 1669390400
transform -1 0 78848 0 1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1669390400
transform 1 0 76720 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1461_
timestamp 1669390400
transform -1 0 96656 0 -1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1669390400
transform 1 0 95536 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1463_
timestamp 1669390400
transform 1 0 94976 0 -1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_
timestamp 1669390400
transform 1 0 94080 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1465_
timestamp 1669390400
transform -1 0 74144 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1466_
timestamp 1669390400
transform -1 0 92624 0 1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1669390400
transform 1 0 91504 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1468_
timestamp 1669390400
transform 1 0 94528 0 -1 70560
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1469_
timestamp 1669390400
transform 1 0 94640 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1470_
timestamp 1669390400
transform 1 0 71904 0 1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1669390400
transform -1 0 71008 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1472_
timestamp 1669390400
transform -1 0 90832 0 -1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1473_
timestamp 1669390400
transform -1 0 93744 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1474_
timestamp 1669390400
transform -1 0 72800 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1475_
timestamp 1669390400
transform 1 0 61264 0 1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1476_
timestamp 1669390400
transform 1 0 60144 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1477_
timestamp 1669390400
transform 1 0 70000 0 1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1478_
timestamp 1669390400
transform 1 0 68432 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1479_
timestamp 1669390400
transform 1 0 61488 0 1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1669390400
transform 1 0 60144 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1481_
timestamp 1669390400
transform -1 0 65072 0 1 72128
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1482_
timestamp 1669390400
transform -1 0 62720 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1483_
timestamp 1669390400
transform 1 0 73584 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1484_
timestamp 1669390400
transform 1 0 61264 0 1 67424
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1485_
timestamp 1669390400
transform -1 0 60816 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1486_
timestamp 1669390400
transform 1 0 61936 0 -1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1669390400
transform -1 0 61712 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1488_
timestamp 1669390400
transform -1 0 77616 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1489_
timestamp 1669390400
transform 1 0 76160 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1490_
timestamp 1669390400
transform 1 0 61376 0 1 65856
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1491_
timestamp 1669390400
transform 1 0 60144 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1492_
timestamp 1669390400
transform 1 0 73360 0 -1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1493_
timestamp 1669390400
transform 1 0 75600 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1494_
timestamp 1669390400
transform 1 0 94976 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1495_
timestamp 1669390400
transform 1 0 94080 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1496_
timestamp 1669390400
transform 1 0 76496 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1497_
timestamp 1669390400
transform 1 0 77168 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1498_
timestamp 1669390400
transform -1 0 92288 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1499_
timestamp 1669390400
transform -1 0 93296 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1500_
timestamp 1669390400
transform 1 0 94976 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1501_
timestamp 1669390400
transform 1 0 94080 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1502_
timestamp 1669390400
transform -1 0 75040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1503_
timestamp 1669390400
transform 1 0 84000 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1504_
timestamp 1669390400
transform -1 0 84336 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1505_
timestamp 1669390400
transform 1 0 89600 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1506_
timestamp 1669390400
transform 1 0 89600 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1507_
timestamp 1669390400
transform 1 0 68992 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1508_
timestamp 1669390400
transform -1 0 68208 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1509_
timestamp 1669390400
transform 1 0 86464 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1669390400
transform -1 0 88144 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1511_
timestamp 1669390400
transform -1 0 72800 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1512_
timestamp 1669390400
transform 1 0 57792 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1513_
timestamp 1669390400
transform -1 0 56112 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1514_
timestamp 1669390400
transform 1 0 67088 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1515_
timestamp 1669390400
transform -1 0 67200 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1516_
timestamp 1669390400
transform 1 0 51744 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1517_
timestamp 1669390400
transform -1 0 51856 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1518_
timestamp 1669390400
transform 1 0 55216 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1519_
timestamp 1669390400
transform -1 0 54992 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1520_
timestamp 1669390400
transform 1 0 73696 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1521_
timestamp 1669390400
transform 1 0 50848 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1522_
timestamp 1669390400
transform 1 0 48720 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1523_
timestamp 1669390400
transform 1 0 53312 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1524_
timestamp 1669390400
transform -1 0 51520 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1525_
timestamp 1669390400
transform -1 0 76048 0 1 68992
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1526_
timestamp 1669390400
transform 1 0 75040 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1527_
timestamp 1669390400
transform 1 0 51072 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1528_
timestamp 1669390400
transform -1 0 50848 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1529_
timestamp 1669390400
transform 1 0 73248 0 -1 65856
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1530_
timestamp 1669390400
transform 1 0 76608 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1531_
timestamp 1669390400
transform 1 0 82992 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1532_
timestamp 1669390400
transform -1 0 78624 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1533_
timestamp 1669390400
transform 1 0 77616 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1534_
timestamp 1669390400
transform 1 0 85680 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1535_
timestamp 1669390400
transform -1 0 84560 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1536_
timestamp 1669390400
transform -1 0 81760 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1537_
timestamp 1669390400
transform 1 0 78960 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1538_
timestamp 1669390400
transform 1 0 79744 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1539_
timestamp 1669390400
transform 1 0 83440 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1540_
timestamp 1669390400
transform 1 0 86240 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1541_
timestamp 1669390400
transform -1 0 85680 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1542_
timestamp 1669390400
transform -1 0 75040 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1543_
timestamp 1669390400
transform -1 0 89712 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1544_
timestamp 1669390400
transform -1 0 88368 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1545_
timestamp 1669390400
transform 1 0 83104 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1546_
timestamp 1669390400
transform 1 0 88592 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1547_
timestamp 1669390400
transform -1 0 84672 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1548_
timestamp 1669390400
transform -1 0 91168 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1549_
timestamp 1669390400
transform -1 0 88032 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1550_
timestamp 1669390400
transform -1 0 72352 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1551_
timestamp 1669390400
transform 1 0 67424 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1552_
timestamp 1669390400
transform -1 0 75152 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1553_
timestamp 1669390400
transform -1 0 68768 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1554_
timestamp 1669390400
transform -1 0 67984 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1555_
timestamp 1669390400
transform -1 0 90496 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1556_
timestamp 1669390400
transform 1 0 90048 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1557_
timestamp 1669390400
transform -1 0 53088 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1558_
timestamp 1669390400
transform 1 0 51744 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1559_
timestamp 1669390400
transform -1 0 52416 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1560_
timestamp 1669390400
transform -1 0 70448 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1669390400
transform -1 0 68768 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1562_
timestamp 1669390400
transform -1 0 50624 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1563_
timestamp 1669390400
transform 1 0 50960 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1564_
timestamp 1669390400
transform -1 0 50400 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1565_
timestamp 1669390400
transform 1 0 75376 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1566_
timestamp 1669390400
transform -1 0 55552 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1669390400
transform -1 0 54320 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1568_
timestamp 1669390400
transform -1 0 52752 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1569_
timestamp 1669390400
transform -1 0 53424 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1570_
timestamp 1669390400
transform 1 0 49056 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1571_
timestamp 1669390400
transform -1 0 52640 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1572_
timestamp 1669390400
transform -1 0 51968 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1573_
timestamp 1669390400
transform -1 0 76160 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1574_
timestamp 1669390400
transform -1 0 77056 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1575_
timestamp 1669390400
transform -1 0 53872 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1576_
timestamp 1669390400
transform -1 0 51184 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1577_
timestamp 1669390400
transform 1 0 72576 0 1 64288
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1578_
timestamp 1669390400
transform 1 0 75040 0 1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1669390400
transform -1 0 83552 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1580_
timestamp 1669390400
transform 1 0 71792 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1669390400
transform 1 0 73360 0 -1 81536
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1669390400
transform -1 0 82656 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1583_
timestamp 1669390400
transform -1 0 81760 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1584_
timestamp 1669390400
transform -1 0 76496 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1585_
timestamp 1669390400
transform -1 0 75488 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1586_
timestamp 1669390400
transform -1 0 74816 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1587_
timestamp 1669390400
transform -1 0 83888 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1588_
timestamp 1669390400
transform 1 0 82320 0 1 86240
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1589_
timestamp 1669390400
transform -1 0 81648 0 1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1590_
timestamp 1669390400
transform -1 0 71904 0 -1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1591_
timestamp 1669390400
transform -1 0 83440 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1592_
timestamp 1669390400
transform 1 0 80192 0 -1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1669390400
transform -1 0 84336 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1594_
timestamp 1669390400
transform -1 0 82096 0 1 86240
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1595_
timestamp 1669390400
transform 1 0 83440 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1596_
timestamp 1669390400
transform 1 0 83440 0 1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1669390400
transform -1 0 85232 0 -1 84672
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1598_
timestamp 1669390400
transform -1 0 69552 0 -1 78400
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1599_
timestamp 1669390400
transform 1 0 67648 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1600_
timestamp 1669390400
transform -1 0 72800 0 -1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1669390400
transform -1 0 69776 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1602_
timestamp 1669390400
transform -1 0 70336 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1603_
timestamp 1669390400
transform -1 0 83216 0 1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1669390400
transform 1 0 80192 0 -1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1605_
timestamp 1669390400
transform 1 0 50512 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1606_
timestamp 1669390400
transform -1 0 53424 0 -1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1607_
timestamp 1669390400
transform -1 0 52640 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1608_
timestamp 1669390400
transform -1 0 70560 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1669390400
transform 1 0 67872 0 1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1669390400
transform 1 0 49504 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1611_
timestamp 1669390400
transform -1 0 53872 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1612_
timestamp 1669390400
transform -1 0 50512 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1613_
timestamp 1669390400
transform 1 0 70336 0 -1 79968
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1614_
timestamp 1669390400
transform -1 0 57344 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1615_
timestamp 1669390400
transform -1 0 55552 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1616_
timestamp 1669390400
transform 1 0 50288 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1617_
timestamp 1669390400
transform -1 0 53872 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1618_
timestamp 1669390400
transform -1 0 51296 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1619_
timestamp 1669390400
transform -1 0 54880 0 -1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1620_
timestamp 1669390400
transform -1 0 54656 0 1 83104
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1621_
timestamp 1669390400
transform 1 0 75824 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1669390400
transform 1 0 79520 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1623_
timestamp 1669390400
transform -1 0 56336 0 -1 81536
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1624_
timestamp 1669390400
transform -1 0 55664 0 -1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1669390400
transform -1 0 83664 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1626_
timestamp 1669390400
transform 1 0 84112 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1669390400
transform -1 0 83552 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1628_
timestamp 1669390400
transform 1 0 75376 0 1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1669390400
transform -1 0 78512 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1630_
timestamp 1669390400
transform -1 0 77728 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1669390400
transform 1 0 82880 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1669390400
transform 1 0 85120 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1633_
timestamp 1669390400
transform -1 0 84560 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1669390400
transform 1 0 85904 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1669390400
transform 1 0 86800 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1636_
timestamp 1669390400
transform -1 0 82880 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1669390400
transform -1 0 82544 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1638_
timestamp 1669390400
transform -1 0 81760 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1639_
timestamp 1669390400
transform 1 0 84112 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1640_
timestamp 1669390400
transform -1 0 89712 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1641_
timestamp 1669390400
transform -1 0 65968 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1642_
timestamp 1669390400
transform 1 0 64288 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1643_
timestamp 1669390400
transform -1 0 72464 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1669390400
transform -1 0 67536 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1645_
timestamp 1669390400
transform -1 0 66752 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1669390400
transform -1 0 83104 0 1 79968
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1647_
timestamp 1669390400
transform -1 0 81984 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1648_
timestamp 1669390400
transform -1 0 52640 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1669390400
transform -1 0 54656 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1650_
timestamp 1669390400
transform -1 0 52416 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1651_
timestamp 1669390400
transform -1 0 65968 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1669390400
transform -1 0 66640 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1653_
timestamp 1669390400
transform -1 0 65856 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1654_
timestamp 1669390400
transform 1 0 51072 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1669390400
transform -1 0 53872 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1656_
timestamp 1669390400
transform -1 0 51856 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1657_
timestamp 1669390400
transform -1 0 56896 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1658_
timestamp 1669390400
transform -1 0 56224 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1659_
timestamp 1669390400
transform 1 0 50512 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1660_
timestamp 1669390400
transform -1 0 55440 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1661_
timestamp 1669390400
transform -1 0 51856 0 1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1662_
timestamp 1669390400
transform -1 0 58688 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1669390400
transform -1 0 55216 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1664_
timestamp 1669390400
transform 1 0 71680 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1669390400
transform 1 0 72576 0 1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1666_
timestamp 1669390400
transform -1 0 58352 0 -1 78400
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1667_
timestamp 1669390400
transform -1 0 57904 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1668_
timestamp 1669390400
transform 1 0 72016 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1669_
timestamp 1669390400
transform 1 0 73696 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1670_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 81200 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1671_
timestamp 1669390400
transform 1 0 77504 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1672_
timestamp 1669390400
transform 1 0 81648 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1673_
timestamp 1669390400
transform 1 0 84672 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1674_
timestamp 1669390400
transform 1 0 81200 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1675_
timestamp 1669390400
transform 1 0 85120 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1676_
timestamp 1669390400
transform 1 0 63952 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1677_
timestamp 1669390400
transform 1 0 82320 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1678_
timestamp 1669390400
transform 1 0 48160 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1679_
timestamp 1669390400
transform 1 0 63840 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1680_
timestamp 1669390400
transform 1 0 48160 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1681_
timestamp 1669390400
transform 1 0 49392 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1682_
timestamp 1669390400
transform 1 0 48160 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1683_
timestamp 1669390400
transform 1 0 48608 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1684_
timestamp 1669390400
transform 1 0 49392 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1685_
timestamp 1669390400
transform -1 0 98000 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1686_
timestamp 1669390400
transform 1 0 76944 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1687_
timestamp 1669390400
transform -1 0 89824 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1688_
timestamp 1669390400
transform -1 0 98000 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1689_
timestamp 1669390400
transform 1 0 81200 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1690_
timestamp 1669390400
transform 1 0 84672 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1691_
timestamp 1669390400
transform 1 0 67200 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1692_
timestamp 1669390400
transform 1 0 82320 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1693_
timestamp 1669390400
transform 1 0 58464 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1694_
timestamp 1669390400
transform 1 0 66192 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1695_
timestamp 1669390400
transform 1 0 57344 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1696_
timestamp 1669390400
transform 1 0 58688 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1697_
timestamp 1669390400
transform 1 0 48832 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1698_
timestamp 1669390400
transform 1 0 55104 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1699_
timestamp 1669390400
transform 1 0 73472 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1700_
timestamp 1669390400
transform 1 0 49840 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1701_
timestamp 1669390400
transform 1 0 94528 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1702_
timestamp 1669390400
transform 1 0 78288 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1703_
timestamp 1669390400
transform -1 0 92624 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1704_
timestamp 1669390400
transform -1 0 98000 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1705_
timestamp 1669390400
transform 1 0 82096 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1706_
timestamp 1669390400
transform -1 0 92400 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1707_
timestamp 1669390400
transform 1 0 69552 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1708_
timestamp 1669390400
transform 1 0 85120 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1709_
timestamp 1669390400
transform 1 0 60816 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1710_
timestamp 1669390400
transform 1 0 70672 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1711_
timestamp 1669390400
transform 1 0 61264 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1712_
timestamp 1669390400
transform -1 0 65184 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1713_
timestamp 1669390400
transform -1 0 65296 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1714_
timestamp 1669390400
transform 1 0 61936 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1715_
timestamp 1669390400
transform 1 0 69328 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1716_
timestamp 1669390400
transform 1 0 62944 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1717_
timestamp 1669390400
transform -1 0 98000 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1718_
timestamp 1669390400
transform 1 0 78848 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1719_
timestamp 1669390400
transform 1 0 93408 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1720_
timestamp 1669390400
transform -1 0 97888 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1721_
timestamp 1669390400
transform 1 0 94752 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1722_
timestamp 1669390400
transform -1 0 94304 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1723_
timestamp 1669390400
transform 1 0 68544 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1724_
timestamp 1669390400
transform -1 0 97888 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1725_
timestamp 1669390400
transform -1 0 64512 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1726_
timestamp 1669390400
transform 1 0 70896 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1727_
timestamp 1669390400
transform 1 0 61264 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1728_
timestamp 1669390400
transform -1 0 65968 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1729_
timestamp 1669390400
transform 1 0 61264 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1730_
timestamp 1669390400
transform 1 0 61712 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1731_
timestamp 1669390400
transform 1 0 75264 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1732_
timestamp 1669390400
transform 1 0 61600 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1733_
timestamp 1669390400
transform 1 0 93408 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1734_
timestamp 1669390400
transform 1 0 79632 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1735_
timestamp 1669390400
transform 1 0 94080 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1736_
timestamp 1669390400
transform 1 0 93408 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1737_
timestamp 1669390400
transform 1 0 93408 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1738_
timestamp 1669390400
transform 1 0 93744 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1739_
timestamp 1669390400
transform 1 0 65520 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1740_
timestamp 1669390400
transform 1 0 93408 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1741_
timestamp 1669390400
transform 1 0 53648 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1742_
timestamp 1669390400
transform 1 0 66192 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1743_
timestamp 1669390400
transform 1 0 53536 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1744_
timestamp 1669390400
transform 1 0 54992 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1745_
timestamp 1669390400
transform 1 0 53424 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1746_
timestamp 1669390400
transform 1 0 53648 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1747_
timestamp 1669390400
transform 1 0 77392 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1748_
timestamp 1669390400
transform 1 0 53536 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1749_
timestamp 1669390400
transform 1 0 94752 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1750_
timestamp 1669390400
transform 1 0 77504 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1751_
timestamp 1669390400
transform -1 0 96320 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1752_
timestamp 1669390400
transform -1 0 98000 0 1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1753_
timestamp 1669390400
transform 1 0 87696 0 1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1754_
timestamp 1669390400
transform 1 0 89376 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1755_
timestamp 1669390400
transform 1 0 67984 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1756_
timestamp 1669390400
transform 1 0 87472 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1757_
timestamp 1669390400
transform 1 0 54880 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1758_
timestamp 1669390400
transform 1 0 66864 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1759_
timestamp 1669390400
transform 1 0 53648 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1760_
timestamp 1669390400
transform 1 0 56896 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1761_
timestamp 1669390400
transform 1 0 48608 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1762_
timestamp 1669390400
transform 1 0 53424 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1763_
timestamp 1669390400
transform 1 0 78064 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1764_
timestamp 1669390400
transform 1 0 49392 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1765_
timestamp 1669390400
transform 1 0 94752 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1766_
timestamp 1669390400
transform 1 0 77168 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1767_
timestamp 1669390400
transform 1 0 94752 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1768_
timestamp 1669390400
transform 1 0 94752 0 1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1769_
timestamp 1669390400
transform 1 0 90720 0 -1 89376
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1770_
timestamp 1669390400
transform 1 0 94752 0 1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1771_
timestamp 1669390400
transform 1 0 69216 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1772_
timestamp 1669390400
transform -1 0 93744 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1773_
timestamp 1669390400
transform 1 0 56224 0 1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1774_
timestamp 1669390400
transform 1 0 67200 0 -1 87808
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1775_
timestamp 1669390400
transform 1 0 59696 0 -1 87808
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1776_
timestamp 1669390400
transform 1 0 57344 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1777_
timestamp 1669390400
transform 1 0 62720 0 1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1778_
timestamp 1669390400
transform -1 0 64064 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1779_
timestamp 1669390400
transform 1 0 74144 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1780_
timestamp 1669390400
transform -1 0 65744 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1781_
timestamp 1669390400
transform -1 0 94528 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1782_
timestamp 1669390400
transform 1 0 75264 0 -1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1783_
timestamp 1669390400
transform -1 0 94640 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1784_
timestamp 1669390400
transform -1 0 93520 0 -1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1785_
timestamp 1669390400
transform -1 0 88704 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1786_
timestamp 1669390400
transform -1 0 88704 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1787_
timestamp 1669390400
transform 1 0 67984 0 -1 89376
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1788_
timestamp 1669390400
transform 1 0 85120 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1789_
timestamp 1669390400
transform 1 0 50848 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1790_
timestamp 1669390400
transform 1 0 66192 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1791_
timestamp 1669390400
transform 1 0 54208 0 1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1792_
timestamp 1669390400
transform 1 0 50960 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1793_
timestamp 1669390400
transform -1 0 64512 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1794_
timestamp 1669390400
transform 1 0 57344 0 -1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1795_
timestamp 1669390400
transform 1 0 74368 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1796_
timestamp 1669390400
transform 1 0 60368 0 -1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1797_
timestamp 1669390400
transform 1 0 90944 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1798_
timestamp 1669390400
transform 1 0 73808 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1799_
timestamp 1669390400
transform -1 0 91056 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1800_
timestamp 1669390400
transform -1 0 96320 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1801_
timestamp 1669390400
transform 1 0 78064 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1802_
timestamp 1669390400
transform 1 0 81200 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1803_
timestamp 1669390400
transform 1 0 66528 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1804_
timestamp 1669390400
transform 1 0 78624 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1805_
timestamp 1669390400
transform -1 0 60592 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1806_
timestamp 1669390400
transform 1 0 65296 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1807_
timestamp 1669390400
transform 1 0 53648 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1808_
timestamp 1669390400
transform 1 0 55888 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1809_
timestamp 1669390400
transform 1 0 49392 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1810_
timestamp 1669390400
transform 1 0 53872 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1811_
timestamp 1669390400
transform 1 0 73360 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1812_
timestamp 1669390400
transform 1 0 49616 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1813_
timestamp 1669390400
transform 1 0 89488 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1814_
timestamp 1669390400
transform -1 0 76944 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1815_
timestamp 1669390400
transform 1 0 89040 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1816_
timestamp 1669390400
transform -1 0 88704 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1817_
timestamp 1669390400
transform 1 0 89152 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1818_
timestamp 1669390400
transform -1 0 88144 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1819_
timestamp 1669390400
transform 1 0 66752 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1820_
timestamp 1669390400
transform 1 0 81424 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1821_
timestamp 1669390400
transform 1 0 55216 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1822_
timestamp 1669390400
transform 1 0 66640 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1823_
timestamp 1669390400
transform 1 0 49616 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1824_
timestamp 1669390400
transform 1 0 55664 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1825_
timestamp 1669390400
transform 1 0 49168 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1826_
timestamp 1669390400
transform 1 0 51632 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1827_
timestamp 1669390400
transform 1 0 71792 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1828_
timestamp 1669390400
transform 1 0 49616 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1829_
timestamp 1669390400
transform 1 0 89152 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1830_
timestamp 1669390400
transform 1 0 77504 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1831_
timestamp 1669390400
transform -1 0 90944 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1832_
timestamp 1669390400
transform -1 0 92400 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1833_
timestamp 1669390400
transform 1 0 88816 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1834_
timestamp 1669390400
transform -1 0 88368 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1835_
timestamp 1669390400
transform 1 0 66416 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1836_
timestamp 1669390400
transform -1 0 91616 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1837_
timestamp 1669390400
transform 1 0 61488 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1838_
timestamp 1669390400
transform 1 0 67088 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1839_
timestamp 1669390400
transform 1 0 60480 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1840_
timestamp 1669390400
transform 1 0 61264 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1841_
timestamp 1669390400
transform 1 0 61264 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1842_
timestamp 1669390400
transform 1 0 59360 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1843_
timestamp 1669390400
transform 1 0 73472 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1844_
timestamp 1669390400
transform -1 0 64512 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1845_
timestamp 1669390400
transform 1 0 94528 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1846_
timestamp 1669390400
transform 1 0 77392 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1847_
timestamp 1669390400
transform -1 0 98000 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1848_
timestamp 1669390400
transform -1 0 97328 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1849_
timestamp 1669390400
transform -1 0 94080 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1850_
timestamp 1669390400
transform -1 0 96656 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1851_
timestamp 1669390400
transform 1 0 69328 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1852_
timestamp 1669390400
transform -1 0 92624 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1853_
timestamp 1669390400
transform 1 0 60368 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1854_
timestamp 1669390400
transform 1 0 67984 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1855_
timestamp 1669390400
transform 1 0 61264 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1856_
timestamp 1669390400
transform 1 0 61264 0 -1 73696
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1857_
timestamp 1669390400
transform 1 0 59584 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1858_
timestamp 1669390400
transform 1 0 60368 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1859_
timestamp 1669390400
transform 1 0 77168 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1860_
timestamp 1669390400
transform 1 0 59808 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1861_
timestamp 1669390400
transform 1 0 94192 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1862_
timestamp 1669390400
transform -1 0 79072 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1863_
timestamp 1669390400
transform -1 0 92624 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1864_
timestamp 1669390400
transform 1 0 94416 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1865_
timestamp 1669390400
transform 1 0 82992 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1866_
timestamp 1669390400
transform 1 0 89152 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1867_
timestamp 1669390400
transform 1 0 65520 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1868_
timestamp 1669390400
transform 1 0 85568 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1869_
timestamp 1669390400
transform 1 0 54320 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1870_
timestamp 1669390400
transform 1 0 65520 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1871_
timestamp 1669390400
transform 1 0 49616 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1872_
timestamp 1669390400
transform 1 0 53648 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1873_
timestamp 1669390400
transform 1 0 49392 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1874_
timestamp 1669390400
transform 1 0 49840 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1875_
timestamp 1669390400
transform -1 0 77168 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1876_
timestamp 1669390400
transform 1 0 49616 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1877_
timestamp 1669390400
transform 1 0 82992 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1878_
timestamp 1669390400
transform 1 0 78400 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1879_
timestamp 1669390400
transform 1 0 85120 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1880_
timestamp 1669390400
transform 1 0 87696 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1881_
timestamp 1669390400
transform 1 0 85120 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1882_
timestamp 1669390400
transform 1 0 87136 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1883_
timestamp 1669390400
transform 1 0 65968 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1884_
timestamp 1669390400
transform -1 0 91840 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1885_
timestamp 1669390400
transform 1 0 48720 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1886_
timestamp 1669390400
transform 1 0 66416 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1887_
timestamp 1669390400
transform 1 0 48608 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1888_
timestamp 1669390400
transform 1 0 53424 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1889_
timestamp 1669390400
transform 1 0 49392 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1890_
timestamp 1669390400
transform 1 0 49392 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1891_
timestamp 1669390400
transform 1 0 73472 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1892_
timestamp 1669390400
transform 1 0 49168 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1893_
timestamp 1669390400
transform 1 0 78624 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1894_
timestamp 1669390400
transform 1 0 73248 0 -1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1895_
timestamp 1669390400
transform 1 0 79968 0 1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1896_
timestamp 1669390400
transform 1 0 81200 0 -1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1897_
timestamp 1669390400
transform -1 0 84448 0 -1 86240
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1898_
timestamp 1669390400
transform 1 0 81760 0 -1 83104
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1899_
timestamp 1669390400
transform 1 0 65520 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1900_
timestamp 1669390400
transform 1 0 81200 0 -1 84672
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1901_
timestamp 1669390400
transform 1 0 49280 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1902_
timestamp 1669390400
transform -1 0 69440 0 -1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1903_
timestamp 1669390400
transform 1 0 49392 0 -1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1904_
timestamp 1669390400
transform 1 0 53312 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1905_
timestamp 1669390400
transform 1 0 49616 0 1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1906_
timestamp 1669390400
transform 1 0 51520 0 -1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1907_
timestamp 1669390400
transform 1 0 77504 0 -1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1908_
timestamp 1669390400
transform 1 0 53984 0 1 81536
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1909_
timestamp 1669390400
transform 1 0 81648 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1910_
timestamp 1669390400
transform 1 0 73696 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1911_
timestamp 1669390400
transform 1 0 83328 0 -1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1912_
timestamp 1669390400
transform -1 0 88368 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1913_
timestamp 1669390400
transform 1 0 78848 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1914_
timestamp 1669390400
transform -1 0 88592 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1915_
timestamp 1669390400
transform 1 0 63616 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1916_
timestamp 1669390400
transform 1 0 81200 0 -1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1917_
timestamp 1669390400
transform 1 0 49840 0 -1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1918_
timestamp 1669390400
transform 1 0 64176 0 1 78400
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1919_
timestamp 1669390400
transform 1 0 49616 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1920_
timestamp 1669390400
transform 1 0 53648 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1921_
timestamp 1669390400
transform 1 0 49616 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1922_
timestamp 1669390400
transform 1 0 54208 0 1 76832
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1923_
timestamp 1669390400
transform 1 0 71456 0 1 79968
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1924_
timestamp 1669390400
transform 1 0 57120 0 1 75264
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1925_
timestamp 1669390400
transform 1 0 72800 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 78960 0 -1 61152
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1669390400
transform -1 0 62944 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1669390400
transform 1 0 89152 0 -1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1669390400
transform -1 0 62944 0 -1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1669390400
transform 1 0 87024 0 1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1669390400
transform -1 0 56672 0 -1 56448
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1669390400
transform 1 0 58800 0 -1 58016
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1669390400
transform -1 0 67424 0 1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1669390400
transform -1 0 68768 0 1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1669390400
transform -1 0 70896 0 -1 65856
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1669390400
transform -1 0 66864 0 1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1669390400
transform -1 0 55552 0 -1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1669390400
transform 1 0 51296 0 -1 70560
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1669390400
transform 1 0 51296 0 -1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1669390400
transform 1 0 51296 0 -1 83104
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1669390400
transform 1 0 58464 0 -1 84672
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1669390400
transform -1 0 68096 0 1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1669390400
transform 1 0 65856 0 -1 86240
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1669390400
transform 1 0 69216 0 1 78400
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1669390400
transform 1 0 63168 0 1 73696
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1669390400
transform 1 0 69216 0 1 70560
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1669390400
transform -1 0 82768 0 1 67424
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1669390400
transform -1 0 84224 0 1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1669390400
transform -1 0 82768 0 1 78400
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1669390400
transform -1 0 82768 0 1 84672
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1669390400
transform 1 0 85120 0 1 81536
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1669390400
transform -1 0 92624 0 1 79968
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1669390400
transform -1 0 94752 0 -1 87808
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1669390400
transform 1 0 91056 0 -1 83104
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1669390400
transform 1 0 91056 0 -1 76832
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1669390400
transform 1 0 89712 0 -1 72128
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1669390400
transform 1 0 91056 0 -1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1669390400
transform -1 0 96656 0 -1 61152
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_28_clk
timestamp 1669390400
transform -1 0 94752 0 -1 67424
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_clk
timestamp 1669390400
transform -1 0 88704 0 -1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_clk
timestamp 1669390400
transform 1 0 81536 0 -1 56448
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_clk
timestamp 1669390400
transform -1 0 92512 0 1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_clk
timestamp 1669390400
transform 1 0 91056 0 -1 56448
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_clk
timestamp 1669390400
transform 1 0 91056 0 -1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_clk
timestamp 1669390400
transform 1 0 89824 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_clk
timestamp 1669390400
transform 1 0 91056 0 -1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_clk
timestamp 1669390400
transform -1 0 96656 0 -1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_clk
timestamp 1669390400
transform -1 0 95872 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_39_clk
timestamp 1669390400
transform 1 0 83104 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_40_clk
timestamp 1669390400
transform -1 0 86800 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_41_clk
timestamp 1669390400
transform -1 0 80640 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_42_clk
timestamp 1669390400
transform -1 0 84672 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_43_clk
timestamp 1669390400
transform 1 0 77952 0 1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_44_clk
timestamp 1669390400
transform 1 0 69440 0 1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_45_clk
timestamp 1669390400
transform -1 0 68768 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_46_clk
timestamp 1669390400
transform 1 0 69216 0 1 42336
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_47_clk
timestamp 1669390400
transform 1 0 66864 0 -1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_48_clk
timestamp 1669390400
transform 1 0 62160 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_50_clk
timestamp 1669390400
transform 1 0 55216 0 1 34496
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_51_clk
timestamp 1669390400
transform -1 0 55776 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_52_clk
timestamp 1669390400
transform 1 0 53312 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1669390400
transform 1 0 1680 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1669390400
transform 1 0 1680 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1669390400
transform 1 0 1680 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 1 87808
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1669390400
transform 1 0 6496 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1669390400
transform 1 0 18928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1669390400
transform 1 0 31360 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1669390400
transform 1 0 44800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1669390400
transform 1 0 56560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1669390400
transform 1 0 68656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1669390400
transform 1 0 81088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1669390400
transform -1 0 94192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1669390400
transform -1 0 95424 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output14 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8064 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output15
timestamp 1669390400
transform -1 0 20496 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output16
timestamp 1669390400
transform -1 0 32592 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output17
timestamp 1669390400
transform -1 0 46368 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18
timestamp 1669390400
transform -1 0 58128 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 70224 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform -1 0 82656 0 1 95648
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform 1 0 93520 0 1 95648
box -86 -86 1654 870
<< labels >>
flabel metal3 s 0 12432 800 12544 0 FreeSans 448 0 0 0 address[0]
port 0 nsew signal input
flabel metal3 s 0 37408 800 37520 0 FreeSans 448 0 0 0 address[1]
port 1 nsew signal input
flabel metal3 s 0 62384 800 62496 0 FreeSans 448 0 0 0 address[2]
port 2 nsew signal input
flabel metal3 s 0 87360 800 87472 0 FreeSans 448 0 0 0 address[3]
port 3 nsew signal input
flabel metal3 s 99200 74928 100000 75040 0 FreeSans 448 0 0 0 clk
port 4 nsew signal input
flabel metal2 s 6384 0 6496 800 0 FreeSans 448 90 0 0 data_in[0]
port 5 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 data_in[1]
port 6 nsew signal input
flabel metal2 s 31248 0 31360 800 0 FreeSans 448 90 0 0 data_in[2]
port 7 nsew signal input
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 data_in[3]
port 8 nsew signal input
flabel metal2 s 56112 0 56224 800 0 FreeSans 448 90 0 0 data_in[4]
port 9 nsew signal input
flabel metal2 s 68544 0 68656 800 0 FreeSans 448 90 0 0 data_in[5]
port 10 nsew signal input
flabel metal2 s 80976 0 81088 800 0 FreeSans 448 90 0 0 data_in[6]
port 11 nsew signal input
flabel metal2 s 93408 0 93520 800 0 FreeSans 448 90 0 0 data_in[7]
port 12 nsew signal input
flabel metal2 s 6384 99200 6496 100000 0 FreeSans 448 90 0 0 data_out[0]
port 13 nsew signal tristate
flabel metal2 s 18816 99200 18928 100000 0 FreeSans 448 90 0 0 data_out[1]
port 14 nsew signal tristate
flabel metal2 s 31248 99200 31360 100000 0 FreeSans 448 90 0 0 data_out[2]
port 15 nsew signal tristate
flabel metal2 s 43680 99200 43792 100000 0 FreeSans 448 90 0 0 data_out[3]
port 16 nsew signal tristate
flabel metal2 s 56112 99200 56224 100000 0 FreeSans 448 90 0 0 data_out[4]
port 17 nsew signal tristate
flabel metal2 s 68544 99200 68656 100000 0 FreeSans 448 90 0 0 data_out[5]
port 18 nsew signal tristate
flabel metal2 s 80976 99200 81088 100000 0 FreeSans 448 90 0 0 data_out[6]
port 19 nsew signal tristate
flabel metal2 s 93408 99200 93520 100000 0 FreeSans 448 90 0 0 data_out[7]
port 20 nsew signal tristate
flabel metal3 s 99200 24976 100000 25088 0 FreeSans 448 0 0 0 rd_wr
port 21 nsew signal input
flabel metal4 s 4448 3076 4768 96492 0 FreeSans 1280 90 0 0 vdd
port 22 nsew power bidirectional
flabel metal4 s 35168 3076 35488 96492 0 FreeSans 1280 90 0 0 vdd
port 22 nsew power bidirectional
flabel metal4 s 65888 3076 66208 96492 0 FreeSans 1280 90 0 0 vdd
port 22 nsew power bidirectional
flabel metal4 s 96608 3076 96928 96492 0 FreeSans 1280 90 0 0 vdd
port 22 nsew power bidirectional
flabel metal4 s 19808 3076 20128 96492 0 FreeSans 1280 90 0 0 vss
port 23 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 96492 0 FreeSans 1280 90 0 0 vss
port 23 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 96492 0 FreeSans 1280 90 0 0 vss
port 23 nsew ground bidirectional
rlabel metal1 49952 96432 49952 96432 0 vdd
rlabel metal1 49952 95648 49952 95648 0 vss
rlabel metal2 82152 45416 82152 45416 0 _0000_
rlabel metal2 78456 45416 78456 45416 0 _0001_
rlabel metal3 83384 54600 83384 54600 0 _0002_
rlabel metal2 85624 44576 85624 44576 0 _0003_
rlabel metal2 82152 72632 82152 72632 0 _0004_
rlabel metal2 85624 54936 85624 54936 0 _0005_
rlabel metal2 64904 69328 64904 69328 0 _0006_
rlabel metal2 83272 71848 83272 71848 0 _0007_
rlabel metal2 49112 60200 49112 60200 0 _0008_
rlabel metal2 64736 64792 64736 64792 0 _0009_
rlabel metal2 49112 57568 49112 57568 0 _0010_
rlabel metal3 49112 59304 49112 59304 0 _0011_
rlabel metal2 48776 54656 48776 54656 0 _0012_
rlabel metal3 48888 53592 48888 53592 0 _0013_
rlabel metal2 49672 52416 49672 52416 0 _0014_
rlabel metal2 97272 42392 97272 42392 0 _0015_
rlabel metal3 77504 43624 77504 43624 0 _0016_
rlabel metal3 89096 40600 89096 40600 0 _0017_
rlabel metal2 97048 44800 97048 44800 0 _0018_
rlabel metal2 81928 37688 81928 37688 0 _0019_
rlabel metal2 85624 41440 85624 41440 0 _0020_
rlabel metal2 68208 39480 68208 39480 0 _0021_
rlabel metal2 83272 39144 83272 39144 0 _0022_
rlabel metal2 59416 39144 59416 39144 0 _0023_
rlabel metal2 67368 41440 67368 41440 0 _0024_
rlabel metal2 57960 41832 57960 41832 0 _0025_
rlabel metal2 59640 42056 59640 42056 0 _0026_
rlabel metal2 48776 43960 48776 43960 0 _0027_
rlabel metal2 56056 44800 56056 44800 0 _0028_
rlabel metal2 74424 76776 74424 76776 0 _0029_
rlabel metal2 50848 45192 50848 45192 0 _0030_
rlabel metal3 94808 37912 94808 37912 0 _0031_
rlabel metal2 79296 39704 79296 39704 0 _0032_
rlabel metal2 91672 36792 91672 36792 0 _0033_
rlabel metal2 97048 40096 97048 40096 0 _0034_
rlabel metal2 83048 32872 83048 32872 0 _0035_
rlabel metal2 89432 37576 89432 37576 0 _0036_
rlabel metal2 70504 34048 70504 34048 0 _0037_
rlabel metal3 85288 34776 85288 34776 0 _0038_
rlabel metal3 61208 33208 61208 33208 0 _0039_
rlabel metal2 71624 31892 71624 31892 0 _0040_
rlabel metal3 61432 35000 61432 35000 0 _0041_
rlabel metal2 64232 33600 64232 33600 0 _0042_
rlabel metal2 64344 41384 64344 41384 0 _0043_
rlabel metal3 63448 38920 63448 38920 0 _0044_
rlabel metal2 70280 43960 70280 43960 0 _0045_
rlabel metal3 63336 42840 63336 42840 0 _0046_
rlabel metal2 97104 49112 97104 49112 0 _0047_
rlabel metal2 79800 49756 79800 49756 0 _0048_
rlabel metal2 93464 47488 93464 47488 0 _0049_
rlabel metal3 96320 53144 96320 53144 0 _0050_
rlabel metal3 95928 50008 95928 50008 0 _0051_
rlabel metal2 93296 49896 93296 49896 0 _0052_
rlabel metal2 69608 50344 69608 50344 0 _0053_
rlabel metal2 97160 51800 97160 51800 0 _0054_
rlabel metal2 63560 45304 63560 45304 0 _0055_
rlabel metal2 71904 50008 71904 50008 0 _0056_
rlabel metal2 60984 47488 60984 47488 0 _0057_
rlabel metal2 65016 46704 65016 46704 0 _0058_
rlabel metal2 62272 45976 62272 45976 0 _0059_
rlabel metal3 62944 50456 62944 50456 0 _0060_
rlabel metal3 75544 38920 75544 38920 0 _0061_
rlabel metal3 63952 49784 63952 49784 0 _0062_
rlabel metal2 94416 55384 94416 55384 0 _0063_
rlabel metal2 80584 56000 80584 56000 0 _0064_
rlabel metal3 94080 56952 94080 56952 0 _0065_
rlabel metal3 96040 59976 96040 59976 0 _0066_
rlabel metal3 94864 57736 94864 57736 0 _0067_
rlabel metal2 92568 60704 92568 60704 0 _0068_
rlabel metal2 66472 55216 66472 55216 0 _0069_
rlabel metal2 94248 60816 94248 60816 0 _0070_
rlabel metal2 54600 56896 54600 56896 0 _0071_
rlabel metal2 67704 60368 67704 60368 0 _0072_
rlabel metal2 54488 55888 54488 55888 0 _0073_
rlabel metal3 55328 58296 55328 58296 0 _0074_
rlabel metal3 53872 56952 53872 56952 0 _0075_
rlabel metal2 54600 60032 54600 60032 0 _0076_
rlabel metal2 78344 50512 78344 50512 0 _0077_
rlabel metal2 54488 59640 54488 59640 0 _0078_
rlabel metal2 95648 74200 95648 74200 0 _0079_
rlabel metal2 78456 72856 78456 72856 0 _0080_
rlabel metal3 94472 75768 94472 75768 0 _0081_
rlabel metal2 97048 73024 97048 73024 0 _0082_
rlabel metal2 88592 74200 88592 74200 0 _0083_
rlabel metal2 90328 76160 90328 76160 0 _0084_
rlabel metal2 69384 75936 69384 75936 0 _0085_
rlabel metal2 88424 72240 88424 72240 0 _0086_
rlabel metal2 55832 71568 55832 71568 0 _0087_
rlabel metal2 68040 74760 68040 74760 0 _0088_
rlabel metal2 54600 71904 54600 71904 0 _0089_
rlabel metal2 56504 69048 56504 69048 0 _0090_
rlabel metal3 48888 70840 48888 70840 0 _0091_
rlabel metal2 54320 68824 54320 68824 0 _0092_
rlabel metal3 79296 56952 79296 56952 0 _0093_
rlabel metal2 50176 69272 50176 69272 0 _0094_
rlabel metal3 96488 79800 96488 79800 0 _0095_
rlabel metal2 78064 84392 78064 84392 0 _0096_
rlabel metal2 95704 85568 95704 85568 0 _0097_
rlabel metal2 95704 78932 95704 78932 0 _0098_
rlabel metal2 91896 87696 91896 87696 0 _0099_
rlabel metal2 95704 84280 95704 84280 0 _0100_
rlabel metal2 70280 84168 70280 84168 0 _0101_
rlabel metal2 93240 85344 93240 85344 0 _0102_
rlabel metal2 57176 87360 57176 87360 0 _0103_
rlabel metal2 68208 86520 68208 86520 0 _0104_
rlabel metal2 61432 86912 61432 86912 0 _0105_
rlabel metal3 59080 85960 59080 85960 0 _0106_
rlabel metal2 63448 83216 63448 83216 0 _0107_
rlabel metal2 61768 85400 61768 85400 0 _0108_
rlabel metal2 75096 73640 75096 73640 0 _0109_
rlabel metal2 64792 85848 64792 85848 0 _0110_
rlabel metal2 93576 78344 93576 78344 0 _0111_
rlabel metal2 76160 82824 76160 82824 0 _0112_
rlabel metal2 93632 83384 93632 83384 0 _0113_
rlabel metal3 92232 79464 92232 79464 0 _0114_
rlabel metal3 87528 85960 87528 85960 0 _0115_
rlabel metal3 88536 84392 88536 84392 0 _0116_
rlabel metal2 69384 86128 69384 86128 0 _0117_
rlabel metal2 86128 85176 86128 85176 0 _0118_
rlabel metal2 51800 85400 51800 85400 0 _0119_
rlabel metal2 68040 84616 68040 84616 0 _0120_
rlabel metal2 55160 85792 55160 85792 0 _0121_
rlabel metal2 52248 85120 52248 85120 0 _0122_
rlabel metal2 63560 80864 63560 80864 0 _0123_
rlabel metal2 58240 82824 58240 82824 0 _0124_
rlabel metal2 75376 85960 75376 85960 0 _0125_
rlabel metal2 61320 82040 61320 82040 0 _0126_
rlabel metal2 91896 39928 91896 39928 0 _0127_
rlabel metal3 76048 41048 76048 41048 0 _0128_
rlabel metal2 89656 39256 89656 39256 0 _0129_
rlabel metal3 94472 41272 94472 41272 0 _0130_
rlabel metal3 80192 32760 80192 32760 0 _0131_
rlabel metal2 82096 42056 82096 42056 0 _0132_
rlabel metal2 68040 36736 68040 36736 0 _0133_
rlabel metal2 79576 34552 79576 34552 0 _0134_
rlabel metal2 59752 34216 59752 34216 0 _0135_
rlabel metal2 66248 38080 66248 38080 0 _0136_
rlabel metal2 55496 39144 55496 39144 0 _0137_
rlabel metal2 56784 36568 56784 36568 0 _0138_
rlabel metal2 49896 41440 49896 41440 0 _0139_
rlabel metal2 54824 43232 54824 43232 0 _0140_
rlabel metal2 74312 84616 74312 84616 0 _0141_
rlabel metal2 50456 41832 50456 41832 0 _0142_
rlabel metal2 90104 46200 90104 46200 0 _0143_
rlabel metal2 76216 46424 76216 46424 0 _0144_
rlabel metal2 90104 47544 90104 47544 0 _0145_
rlabel metal2 87808 46760 87808 46760 0 _0146_
rlabel metal2 90104 49056 90104 49056 0 _0147_
rlabel metal2 87192 49056 87192 49056 0 _0148_
rlabel metal2 67704 45416 67704 45416 0 _0149_
rlabel metal3 82600 48328 82600 48328 0 _0150_
rlabel metal2 56224 45976 56224 45976 0 _0151_
rlabel metal2 68152 46200 68152 46200 0 _0152_
rlabel metal2 50512 48328 50512 48328 0 _0153_
rlabel metal3 57624 48440 57624 48440 0 _0154_
rlabel metal3 51632 47544 51632 47544 0 _0155_
rlabel metal2 54880 47992 54880 47992 0 _0156_
rlabel metal2 72744 40096 72744 40096 0 _0157_
rlabel metal2 50512 49112 50512 49112 0 _0158_
rlabel metal3 89376 56280 89376 56280 0 _0159_
rlabel metal2 78456 55216 78456 55216 0 _0160_
rlabel metal2 89656 53368 89656 53368 0 _0161_
rlabel metal3 90048 57624 90048 57624 0 _0162_
rlabel metal2 89768 55608 89768 55608 0 _0163_
rlabel metal2 87472 53032 87472 53032 0 _0164_
rlabel metal3 67816 53032 67816 53032 0 _0165_
rlabel metal3 90384 58520 90384 58520 0 _0166_
rlabel metal2 64008 55048 64008 55048 0 _0167_
rlabel metal2 68040 51576 68040 51576 0 _0168_
rlabel metal3 61768 54600 61768 54600 0 _0169_
rlabel metal2 62216 57456 62216 57456 0 _0170_
rlabel metal2 62216 53760 62216 53760 0 _0171_
rlabel metal2 60312 58744 60312 58744 0 _0172_
rlabel metal3 75040 44408 75040 44408 0 _0173_
rlabel metal2 63616 58520 63616 58520 0 _0174_
rlabel metal2 94584 65744 94584 65744 0 _0175_
rlabel metal2 77224 69440 77224 69440 0 _0176_
rlabel metal3 96544 69496 96544 69496 0 _0177_
rlabel metal3 95480 64120 95480 64120 0 _0178_
rlabel metal2 93072 70280 93072 70280 0 _0179_
rlabel metal2 95648 67928 95648 67928 0 _0180_
rlabel metal2 70280 72072 70280 72072 0 _0181_
rlabel metal3 92456 69272 92456 69272 0 _0182_
rlabel metal2 60704 73976 60704 73976 0 _0183_
rlabel metal2 68936 71064 68936 71064 0 _0184_
rlabel metal2 60648 71680 60648 71680 0 _0185_
rlabel metal2 62216 74424 62216 74424 0 _0186_
rlabel metal2 60480 67144 60480 67144 0 _0187_
rlabel metal2 61264 68824 61264 68824 0 _0188_
rlabel metal3 77392 53592 77392 53592 0 _0189_
rlabel metal2 60704 65576 60704 65576 0 _0190_
rlabel metal2 94584 34552 94584 34552 0 _0191_
rlabel metal2 77672 33600 77672 33600 0 _0192_
rlabel metal2 91672 33544 91672 33544 0 _0193_
rlabel metal2 95368 34216 95368 34216 0 _0194_
rlabel metal2 83888 31080 83888 31080 0 _0195_
rlabel metal2 90104 32816 90104 32816 0 _0196_
rlabel metal3 67088 31640 67088 31640 0 _0197_
rlabel metal2 86520 33824 86520 33824 0 _0198_
rlabel metal2 55384 31892 55384 31892 0 _0199_
rlabel metal2 66584 33208 66584 33208 0 _0200_
rlabel metal2 51296 33208 51296 33208 0 _0201_
rlabel metal2 54544 32760 54544 32760 0 _0202_
rlabel metal3 49784 37352 49784 37352 0 _0203_
rlabel metal2 51016 34944 51016 34944 0 _0204_
rlabel metal3 75880 70280 75880 70280 0 _0205_
rlabel metal2 50456 38136 50456 38136 0 _0206_
rlabel metal2 84000 65464 84000 65464 0 _0207_
rlabel metal2 79352 67368 79352 67368 0 _0208_
rlabel metal2 85176 67424 85176 67424 0 _0209_
rlabel metal2 88648 65016 88648 65016 0 _0210_
rlabel metal2 84392 69552 84392 69552 0 _0211_
rlabel metal2 88088 66584 88088 66584 0 _0212_
rlabel metal3 67200 67816 67200 67816 0 _0213_
rlabel metal2 90664 69048 90664 69048 0 _0214_
rlabel metal2 49672 68264 49672 68264 0 _0215_
rlabel metal2 67368 68152 67368 68152 0 _0216_
rlabel metal2 49560 65240 49560 65240 0 _0217_
rlabel metal2 53816 65912 53816 65912 0 _0218_
rlabel metal2 50344 65632 50344 65632 0 _0219_
rlabel metal2 50344 64232 50344 64232 0 _0220_
rlabel metal2 74424 35392 74424 35392 0 _0221_
rlabel metal2 50120 63896 50120 63896 0 _0222_
rlabel metal2 79576 80696 79576 80696 0 _0223_
rlabel metal2 74256 79688 74256 79688 0 _0224_
rlabel metal2 81032 81928 81032 81928 0 _0225_
rlabel metal3 81424 79688 81424 79688 0 _0226_
rlabel metal2 83720 84728 83720 84728 0 _0227_
rlabel metal2 82712 83440 82712 83440 0 _0228_
rlabel metal2 69832 78512 69832 78512 0 _0229_
rlabel metal2 80528 82488 80528 82488 0 _0230_
rlabel metal3 51184 78792 51184 78792 0 _0231_
rlabel metal2 68432 81256 68432 81256 0 _0232_
rlabel metal2 50344 80304 50344 80304 0 _0233_
rlabel metal3 54600 80472 54600 80472 0 _0234_
rlabel metal2 50624 81368 50624 81368 0 _0235_
rlabel metal2 52472 82264 52472 82264 0 _0236_
rlabel metal3 79240 65464 79240 65464 0 _0237_
rlabel metal2 55160 80584 55160 80584 0 _0238_
rlabel metal2 83048 74200 83048 74200 0 _0239_
rlabel metal3 75992 77112 75992 77112 0 _0240_
rlabel metal2 84224 76552 84224 76552 0 _0241_
rlabel metal2 87360 76664 87360 76664 0 _0242_
rlabel metal3 80528 75768 80528 75768 0 _0243_
rlabel metal3 88424 78008 88424 78008 0 _0244_
rlabel metal3 65520 75768 65520 75768 0 _0245_
rlabel metal2 81424 77112 81424 77112 0 _0246_
rlabel metal3 51352 74984 51352 74984 0 _0247_
rlabel metal2 65352 78456 65352 78456 0 _0248_
rlabel metal2 51352 75600 51352 75600 0 _0249_
rlabel metal2 54600 75320 54600 75320 0 _0250_
rlabel metal2 50512 75768 50512 75768 0 _0251_
rlabel metal2 55160 77560 55160 77560 0 _0252_
rlabel metal2 72632 80248 72632 80248 0 _0253_
rlabel metal2 58072 75992 58072 75992 0 _0254_
rlabel metal2 73752 46872 73752 46872 0 _0255_
rlabel metal3 87696 85288 87696 85288 0 _0256_
rlabel metal2 54712 86352 54712 86352 0 _0257_
rlabel metal2 52584 86912 52584 86912 0 _0258_
rlabel metal2 68376 85736 68376 85736 0 _0259_
rlabel metal2 55552 86072 55552 86072 0 _0260_
rlabel metal2 52584 85736 52584 85736 0 _0261_
rlabel metal2 73304 81872 73304 81872 0 _0262_
rlabel metal2 63672 80248 63672 80248 0 _0263_
rlabel metal2 58632 82824 58632 82824 0 _0264_
rlabel metal2 74984 85904 74984 85904 0 _0265_
rlabel metal2 62216 82152 62216 82152 0 _0266_
rlabel metal2 72184 57232 72184 57232 0 _0267_
rlabel metal2 72576 53704 72576 53704 0 _0268_
rlabel metal2 76552 39704 76552 39704 0 _0269_
rlabel metal3 94640 41048 94640 41048 0 _0270_
rlabel metal2 74928 38248 74928 38248 0 _0271_
rlabel metal2 89432 39312 89432 39312 0 _0272_
rlabel metal3 92792 42728 92792 42728 0 _0273_
rlabel metal2 71176 36680 71176 36680 0 _0274_
rlabel metal2 81760 32648 81760 32648 0 _0275_
rlabel metal2 82152 41608 82152 41608 0 _0276_
rlabel metal3 68936 36344 68936 36344 0 _0277_
rlabel metal3 81144 34216 81144 34216 0 _0278_
rlabel metal2 68376 38080 68376 38080 0 _0279_
rlabel metal2 59080 36120 59080 36120 0 _0280_
rlabel metal3 66920 37912 66920 37912 0 _0281_
rlabel metal2 56392 38864 56392 38864 0 _0282_
rlabel metal3 57120 37240 57120 37240 0 _0283_
rlabel metal3 53424 41272 53424 41272 0 _0284_
rlabel metal3 50512 41048 50512 41048 0 _0285_
rlabel metal2 55384 42728 55384 42728 0 _0286_
rlabel metal2 74256 83720 74256 83720 0 _0287_
rlabel metal3 51968 41160 51968 41160 0 _0288_
rlabel metal2 72632 63840 72632 63840 0 _0289_
rlabel metal2 71960 63336 71960 63336 0 _0290_
rlabel metal2 71400 51240 71400 51240 0 _0291_
rlabel metal2 78456 49448 78456 49448 0 _0292_
rlabel metal2 94024 47152 94024 47152 0 _0293_
rlabel via2 76440 63896 76440 63896 0 _0294_
rlabel metal2 71456 61992 71456 61992 0 _0295_
rlabel metal2 75768 49448 75768 49448 0 _0296_
rlabel metal2 75544 47208 75544 47208 0 _0297_
rlabel metal2 89768 46536 89768 46536 0 _0298_
rlabel metal2 76496 46872 76496 46872 0 _0299_
rlabel metal3 74928 46872 74928 46872 0 _0300_
rlabel metal2 90216 50232 90216 50232 0 _0301_
rlabel metal2 90776 50120 90776 50120 0 _0302_
rlabel metal2 83944 49224 83944 49224 0 _0303_
rlabel metal3 88088 49784 88088 49784 0 _0304_
rlabel metal2 89432 50176 89432 50176 0 _0305_
rlabel metal2 92680 49112 92680 49112 0 _0306_
rlabel metal3 86184 49000 86184 49000 0 _0307_
rlabel metal2 55272 48496 55272 48496 0 _0308_
rlabel metal2 68488 47768 68488 47768 0 _0309_
rlabel metal2 55272 47320 55272 47320 0 _0310_
rlabel metal3 69328 47320 69328 47320 0 _0311_
rlabel metal2 83384 48888 83384 48888 0 _0312_
rlabel metal3 56952 48328 56952 48328 0 _0313_
rlabel metal2 58408 48272 58408 48272 0 _0314_
rlabel metal2 68488 46480 68488 46480 0 _0315_
rlabel metal3 54264 48776 54264 48776 0 _0316_
rlabel metal2 53704 47992 53704 47992 0 _0317_
rlabel metal2 54488 47656 54488 47656 0 _0318_
rlabel metal2 58184 48328 58184 48328 0 _0319_
rlabel metal2 53368 48496 53368 48496 0 _0320_
rlabel metal2 53480 48384 53480 48384 0 _0321_
rlabel metal2 55048 49280 55048 49280 0 _0322_
rlabel metal2 73584 40376 73584 40376 0 _0323_
rlabel metal2 54376 49504 54376 49504 0 _0324_
rlabel metal2 70728 54936 70728 54936 0 _0325_
rlabel metal2 91280 54488 91280 54488 0 _0326_
rlabel metal2 88480 56168 88480 56168 0 _0327_
rlabel metal2 71512 56392 71512 56392 0 _0328_
rlabel metal2 93464 57512 93464 57512 0 _0329_
rlabel metal3 89320 56168 89320 56168 0 _0330_
rlabel metal2 79016 55776 79016 55776 0 _0331_
rlabel metal2 78736 53144 78736 53144 0 _0332_
rlabel metal2 89488 53144 89488 53144 0 _0333_
rlabel metal3 88424 54712 88424 54712 0 _0334_
rlabel metal3 72072 53480 72072 53480 0 _0335_
rlabel metal2 88312 57960 88312 57960 0 _0336_
rlabel metal3 90384 54712 90384 54712 0 _0337_
rlabel metal2 93128 56504 93128 56504 0 _0338_
rlabel metal2 87304 54096 87304 54096 0 _0339_
rlabel metal2 68488 52080 68488 52080 0 _0340_
rlabel metal2 68152 52192 68152 52192 0 _0341_
rlabel metal2 69608 53480 69608 53480 0 _0342_
rlabel metal2 68600 53032 68600 53032 0 _0343_
rlabel metal2 88648 57120 88648 57120 0 _0344_
rlabel metal2 62888 53872 62888 53872 0 _0345_
rlabel metal2 64344 54656 64344 54656 0 _0346_
rlabel metal2 70056 53032 70056 53032 0 _0347_
rlabel metal3 61040 54712 61040 54712 0 _0348_
rlabel metal2 62440 55104 62440 55104 0 _0349_
rlabel metal2 66920 57456 66920 57456 0 _0350_
rlabel metal3 64120 58632 64120 58632 0 _0351_
rlabel metal2 61656 53312 61656 53312 0 _0352_
rlabel metal3 62048 53144 62048 53144 0 _0353_
rlabel metal3 63112 58296 63112 58296 0 _0354_
rlabel metal2 76328 44408 76328 44408 0 _0355_
rlabel metal2 65352 58520 65352 58520 0 _0356_
rlabel metal2 73528 71960 73528 71960 0 _0357_
rlabel metal3 92568 66360 92568 66360 0 _0358_
rlabel metal2 95312 63672 95312 63672 0 _0359_
rlabel metal2 77000 68880 77000 68880 0 _0360_
rlabel metal3 95480 70392 95480 70392 0 _0361_
rlabel metal2 94808 63896 94808 63896 0 _0362_
rlabel metal2 91336 71008 91336 71008 0 _0363_
rlabel metal2 92344 72240 92344 72240 0 _0364_
rlabel metal2 94808 70616 94808 70616 0 _0365_
rlabel metal2 72184 71008 72184 71008 0 _0366_
rlabel metal2 93464 69160 93464 69160 0 _0367_
rlabel metal2 71288 69552 71288 69552 0 _0368_
rlabel metal3 60984 74088 60984 74088 0 _0369_
rlabel metal3 69496 69608 69496 69608 0 _0370_
rlabel metal3 61096 72520 61096 72520 0 _0371_
rlabel metal2 64792 72856 64792 72856 0 _0372_
rlabel via2 63560 68600 63560 68600 0 _0373_
rlabel metal3 61096 67704 61096 67704 0 _0374_
rlabel metal3 61880 68600 61880 68600 0 _0375_
rlabel metal2 76328 54264 76328 54264 0 _0376_
rlabel metal3 61040 66248 61040 66248 0 _0377_
rlabel metal2 74256 37464 74256 37464 0 _0378_
rlabel metal2 76384 31864 76384 31864 0 _0379_
rlabel metal2 95256 32928 95256 32928 0 _0380_
rlabel metal3 77056 32760 77056 32760 0 _0381_
rlabel metal3 92568 34216 92568 34216 0 _0382_
rlabel metal3 94808 34328 94808 34328 0 _0383_
rlabel metal2 74312 33264 74312 33264 0 _0384_
rlabel metal2 84224 29624 84224 29624 0 _0385_
rlabel metal2 89880 32032 89880 32032 0 _0386_
rlabel metal3 68656 32312 68656 32312 0 _0387_
rlabel metal2 86744 33208 86744 33208 0 _0388_
rlabel metal3 53480 33432 53480 33432 0 _0389_
rlabel metal3 57008 33096 57008 33096 0 _0390_
rlabel metal2 67368 33936 67368 33936 0 _0391_
rlabel metal2 51688 33600 51688 33600 0 _0392_
rlabel metal3 55160 32536 55160 32536 0 _0393_
rlabel metal2 52920 38920 52920 38920 0 _0394_
rlabel metal3 50064 36680 50064 36680 0 _0395_
rlabel metal2 51352 34832 51352 34832 0 _0396_
rlabel metal2 75544 69608 75544 69608 0 _0397_
rlabel metal2 51016 38808 51016 38808 0 _0398_
rlabel metal2 74760 66976 74760 66976 0 _0399_
rlabel metal3 79352 67032 79352 67032 0 _0400_
rlabel metal3 83776 66136 83776 66136 0 _0401_
rlabel metal2 77784 67200 77784 67200 0 _0402_
rlabel metal2 88760 69048 88760 69048 0 _0403_
rlabel metal2 86184 65856 86184 65856 0 _0404_
rlabel metal3 80696 67144 80696 67144 0 _0405_
rlabel metal2 79856 68600 79856 68600 0 _0406_
rlabel metal3 84672 67256 84672 67256 0 _0407_
rlabel metal3 87248 67144 87248 67144 0 _0408_
rlabel metal3 91224 66136 91224 66136 0 _0409_
rlabel metal3 88704 65464 88704 65464 0 _0410_
rlabel metal3 84000 69160 84000 69160 0 _0411_
rlabel metal2 90328 69832 90328 69832 0 _0412_
rlabel metal2 90888 66752 90888 66752 0 _0413_
rlabel metal2 67592 68432 67592 68432 0 _0414_
rlabel metal2 67704 67872 67704 67872 0 _0415_
rlabel metal2 68600 67592 68600 67592 0 _0416_
rlabel metal2 68488 68600 68488 68600 0 _0417_
rlabel metal2 90104 70168 90104 70168 0 _0418_
rlabel metal2 52584 67648 52584 67648 0 _0419_
rlabel metal2 52304 67032 52304 67032 0 _0420_
rlabel metal2 69944 67256 69944 67256 0 _0421_
rlabel metal2 50120 66584 50120 66584 0 _0422_
rlabel metal2 51688 66584 51688 66584 0 _0423_
rlabel metal2 55832 65856 55832 65856 0 _0424_
rlabel metal3 54600 65576 54600 65576 0 _0425_
rlabel metal3 50792 66024 50792 66024 0 _0426_
rlabel metal2 49224 65912 49224 65912 0 _0427_
rlabel metal2 52080 64680 52080 64680 0 _0428_
rlabel metal2 76776 35616 76776 35616 0 _0429_
rlabel metal3 52192 64680 52192 64680 0 _0430_
rlabel metal3 74704 78680 74704 78680 0 _0431_
rlabel metal3 76552 78680 76552 78680 0 _0432_
rlabel metal3 82208 80248 82208 80248 0 _0433_
rlabel metal2 73248 77896 73248 77896 0 _0434_
rlabel metal2 75320 80864 75320 80864 0 _0435_
rlabel metal3 81032 81144 81032 81144 0 _0436_
rlabel metal3 75376 80584 75376 80584 0 _0437_
rlabel metal2 72912 77112 72912 77112 0 _0438_
rlabel metal3 82376 80584 82376 80584 0 _0439_
rlabel metal2 82824 86016 82824 86016 0 _0440_
rlabel metal2 71400 80472 71400 80472 0 _0441_
rlabel metal2 80360 80248 80360 80248 0 _0442_
rlabel metal2 83776 83272 83776 83272 0 _0443_
rlabel via2 82040 83384 82040 83384 0 _0444_
rlabel metal2 83944 82320 83944 82320 0 _0445_
rlabel metal2 50456 78176 50456 78176 0 _0446_
rlabel metal3 69104 78232 69104 78232 0 _0447_
rlabel metal2 53704 78456 53704 78456 0 _0448_
rlabel metal3 68768 80136 68768 80136 0 _0449_
rlabel metal3 81536 81928 81536 81928 0 _0450_
rlabel metal3 51688 78568 51688 78568 0 _0451_
rlabel metal2 52472 78876 52472 78876 0 _0452_
rlabel metal3 69048 80360 69048 80360 0 _0453_
rlabel metal2 50120 81256 50120 81256 0 _0454_
rlabel metal3 53816 78792 53816 78792 0 _0455_
rlabel metal3 71344 77224 71344 77224 0 _0456_
rlabel metal2 55384 80752 55384 80752 0 _0457_
rlabel metal2 50848 78232 50848 78232 0 _0458_
rlabel metal2 53424 83272 53424 83272 0 _0459_
rlabel metal2 54376 80024 54376 80024 0 _0460_
rlabel metal3 77896 65576 77896 65576 0 _0461_
rlabel metal2 55496 80416 55496 80416 0 _0462_
rlabel metal2 83216 73864 83216 73864 0 _0463_
rlabel metal2 84616 75600 84616 75600 0 _0464_
rlabel metal3 76832 76664 76832 76664 0 _0465_
rlabel metal2 77784 77112 77784 77112 0 _0466_
rlabel metal3 83832 77000 83832 77000 0 _0467_
rlabel metal2 84392 77280 84392 77280 0 _0468_
rlabel metal3 86688 75656 86688 75656 0 _0469_
rlabel metal3 81928 75656 81928 75656 0 _0470_
rlabel metal2 81592 76328 81592 76328 0 _0471_
rlabel metal3 87080 78120 87080 78120 0 _0472_
rlabel metal2 52472 74144 52472 74144 0 _0473_
rlabel metal3 65632 76552 65632 76552 0 _0474_
rlabel metal2 55272 74816 55272 74816 0 _0475_
rlabel metal2 66584 76776 66584 76776 0 _0476_
rlabel metal2 82096 77112 82096 77112 0 _0477_
rlabel metal2 52136 75824 52136 75824 0 _0478_
rlabel metal3 53200 75096 53200 75096 0 _0479_
rlabel metal2 66696 78008 66696 78008 0 _0480_
rlabel metal2 65912 78008 65912 78008 0 _0481_
rlabel metal2 51576 75936 51576 75936 0 _0482_
rlabel metal2 53368 75152 53368 75152 0 _0483_
rlabel metal2 56056 76496 56056 76496 0 _0484_
rlabel metal2 51128 73976 51128 73976 0 _0485_
rlabel metal2 54264 77840 54264 77840 0 _0486_
rlabel metal2 55272 77336 55272 77336 0 _0487_
rlabel metal3 72464 77112 72464 77112 0 _0488_
rlabel metal2 57792 76552 57792 76552 0 _0489_
rlabel metal3 73192 46760 73192 46760 0 _0490_
rlabel metal2 72632 59584 72632 59584 0 _0491_
rlabel metal2 78288 64568 78288 64568 0 _0492_
rlabel metal2 87080 65184 87080 65184 0 _0493_
rlabel metal2 78568 61656 78568 61656 0 _0494_
rlabel metal2 77784 77672 77784 77672 0 _0495_
rlabel metal3 69048 59976 69048 59976 0 _0496_
rlabel metal2 68488 77392 68488 77392 0 _0497_
rlabel metal2 78792 77504 78792 77504 0 _0498_
rlabel metal2 78456 76496 78456 76496 0 _0499_
rlabel metal3 81592 64120 81592 64120 0 _0500_
rlabel metal2 73080 57624 73080 57624 0 _0501_
rlabel metal2 69720 64904 69720 64904 0 _0502_
rlabel metal2 86296 64008 86296 64008 0 _0503_
rlabel metal2 69944 60480 69944 60480 0 _0504_
rlabel metal2 66920 60928 66920 60928 0 _0505_
rlabel metal2 90776 63168 90776 63168 0 _0506_
rlabel metal3 80864 62440 80864 62440 0 _0507_
rlabel metal2 70504 62944 70504 62944 0 _0508_
rlabel metal3 71456 62104 71456 62104 0 _0509_
rlabel metal2 86072 63840 86072 63840 0 _0510_
rlabel metal2 81648 62552 81648 62552 0 _0511_
rlabel metal2 68936 63504 68936 63504 0 _0512_
rlabel metal2 73864 52864 73864 52864 0 _0513_
rlabel metal2 77672 48440 77672 48440 0 _0514_
rlabel metal2 73640 53480 73640 53480 0 _0515_
rlabel metal2 78792 49224 78792 49224 0 _0516_
rlabel metal3 79240 48440 79240 48440 0 _0517_
rlabel metal3 80920 64008 80920 64008 0 _0518_
rlabel metal2 86968 62832 86968 62832 0 _0519_
rlabel via2 71624 75768 71624 75768 0 _0520_
rlabel metal2 72184 76216 72184 76216 0 _0521_
rlabel metal2 86408 59920 86408 59920 0 _0522_
rlabel metal2 80416 59864 80416 59864 0 _0523_
rlabel metal2 72184 60816 72184 60816 0 _0524_
rlabel metal2 70504 60928 70504 60928 0 _0525_
rlabel metal2 79800 62328 79800 62328 0 _0526_
rlabel metal3 81032 63896 81032 63896 0 _0527_
rlabel metal3 86800 69832 86800 69832 0 _0528_
rlabel metal2 85288 63784 85288 63784 0 _0529_
rlabel metal2 90328 62776 90328 62776 0 _0530_
rlabel metal2 86520 63448 86520 63448 0 _0531_
rlabel metal3 86856 47208 86856 47208 0 _0532_
rlabel metal3 85288 63000 85288 63000 0 _0533_
rlabel metal2 85848 61040 85848 61040 0 _0534_
rlabel metal2 85848 62944 85848 62944 0 _0535_
rlabel metal2 88312 66248 88312 66248 0 _0536_
rlabel metal2 71568 78008 71568 78008 0 _0537_
rlabel metal2 87528 72464 87528 72464 0 _0538_
rlabel metal3 86520 62384 86520 62384 0 _0539_
rlabel metal2 88312 61880 88312 61880 0 _0540_
rlabel metal3 88480 64120 88480 64120 0 _0541_
rlabel metal2 86520 62552 86520 62552 0 _0542_
rlabel metal2 87136 52024 87136 52024 0 _0543_
rlabel metal2 86296 62608 86296 62608 0 _0544_
rlabel metal2 69272 61712 69272 61712 0 _0545_
rlabel metal2 71512 59360 71512 59360 0 _0546_
rlabel metal3 84280 57736 84280 57736 0 _0547_
rlabel metal3 85008 62328 85008 62328 0 _0548_
rlabel metal2 86744 76328 86744 76328 0 _0549_
rlabel metal2 83048 64680 83048 64680 0 _0550_
rlabel metal3 88480 62440 88480 62440 0 _0551_
rlabel metal2 87640 63280 87640 63280 0 _0552_
rlabel metal2 82376 50064 82376 50064 0 _0553_
rlabel metal3 83832 62552 83832 62552 0 _0554_
rlabel metal3 63616 62440 63616 62440 0 _0555_
rlabel metal2 86240 59864 86240 59864 0 _0556_
rlabel metal2 85736 61936 85736 61936 0 _0557_
rlabel metal2 67704 78596 67704 78596 0 _0558_
rlabel metal2 69216 67928 69216 67928 0 _0559_
rlabel metal3 68824 66136 68824 66136 0 _0560_
rlabel metal3 68992 64568 68992 64568 0 _0561_
rlabel metal2 68376 64624 68376 64624 0 _0562_
rlabel metal2 67928 63560 67928 63560 0 _0563_
rlabel metal2 58632 61824 58632 61824 0 _0564_
rlabel metal2 68096 63224 68096 63224 0 _0565_
rlabel metal2 55048 52024 55048 52024 0 _0566_
rlabel metal2 70840 52696 70840 52696 0 _0567_
rlabel metal2 70952 52024 70952 52024 0 _0568_
rlabel metal3 69496 64680 69496 64680 0 _0569_
rlabel metal2 67312 60872 67312 60872 0 _0570_
rlabel metal2 67928 59472 67928 59472 0 _0571_
rlabel metal3 68600 61544 68600 61544 0 _0572_
rlabel metal2 67760 61656 67760 61656 0 _0573_
rlabel metal2 58576 76664 58576 76664 0 _0574_
rlabel metal2 59640 64288 59640 64288 0 _0575_
rlabel metal2 58464 64120 58464 64120 0 _0576_
rlabel metal2 59248 63112 59248 63112 0 _0577_
rlabel metal2 60256 61096 60256 61096 0 _0578_
rlabel metal2 59696 62552 59696 62552 0 _0579_
rlabel metal2 64904 60200 64904 60200 0 _0580_
rlabel metal2 60088 62776 60088 62776 0 _0581_
rlabel metal3 60032 77672 60032 77672 0 _0582_
rlabel metal3 58408 64456 58408 64456 0 _0583_
rlabel metal3 72632 61880 72632 61880 0 _0584_
rlabel metal2 72016 62328 72016 62328 0 _0585_
rlabel metal2 57400 62832 57400 62832 0 _0586_
rlabel metal2 57624 63000 57624 63000 0 _0587_
rlabel metal2 57400 50736 57400 50736 0 _0588_
rlabel metal3 57960 63112 57960 63112 0 _0589_
rlabel metal2 62888 61656 62888 61656 0 _0590_
rlabel metal2 61936 62552 61936 62552 0 _0591_
rlabel metal2 60312 76020 60312 76020 0 _0592_
rlabel metal2 58520 63112 58520 63112 0 _0593_
rlabel metal2 54712 63784 54712 63784 0 _0594_
rlabel metal2 58184 63224 58184 63224 0 _0595_
rlabel metal2 55608 53648 55608 53648 0 _0596_
rlabel metal3 56896 62552 56896 62552 0 _0597_
rlabel metal2 62440 61432 62440 61432 0 _0598_
rlabel metal2 58856 62944 58856 62944 0 _0599_
rlabel metal2 82544 46872 82544 46872 0 _0600_
rlabel metal3 71736 61544 71736 61544 0 _0601_
rlabel metal2 73472 57848 73472 57848 0 _0602_
rlabel metal2 75768 57904 75768 57904 0 _0603_
rlabel metal2 73864 56504 73864 56504 0 _0604_
rlabel metal2 73528 58520 73528 58520 0 _0605_
rlabel metal3 70784 55384 70784 55384 0 _0606_
rlabel metal2 77952 44184 77952 44184 0 _0607_
rlabel metal2 81816 45864 81816 45864 0 _0608_
rlabel metal2 77448 45136 77448 45136 0 _0609_
rlabel metal3 83328 74536 83328 74536 0 _0610_
rlabel metal2 84224 53928 84224 53928 0 _0611_
rlabel metal2 85400 44968 85400 44968 0 _0612_
rlabel metal3 83328 75432 83328 75432 0 _0613_
rlabel metal2 68600 56280 68600 56280 0 _0614_
rlabel metal2 81872 71176 81872 71176 0 _0615_
rlabel metal3 84896 54600 84896 54600 0 _0616_
rlabel metal2 67928 78736 67928 78736 0 _0617_
rlabel metal2 66248 70616 66248 70616 0 _0618_
rlabel metal2 85400 71512 85400 71512 0 _0619_
rlabel metal3 50064 78680 50064 78680 0 _0620_
rlabel metal2 50568 58464 50568 58464 0 _0621_
rlabel metal3 48944 60872 48944 60872 0 _0622_
rlabel metal3 65016 65576 65016 65576 0 _0623_
rlabel metal2 50288 67256 50288 67256 0 _0624_
rlabel metal3 49000 58408 49000 58408 0 _0625_
rlabel metal2 47656 59864 47656 59864 0 _0626_
rlabel metal2 51464 55160 51464 55160 0 _0627_
rlabel metal2 53928 54208 53928 54208 0 _0628_
rlabel metal2 48384 54600 48384 54600 0 _0629_
rlabel metal2 47992 53984 47992 53984 0 _0630_
rlabel metal2 49336 53144 49336 53144 0 _0631_
rlabel metal2 98000 40600 98000 40600 0 _0632_
rlabel metal3 68432 58408 68432 58408 0 _0633_
rlabel metal2 73528 51800 73528 51800 0 _0634_
rlabel metal2 78008 42672 78008 42672 0 _0635_
rlabel metal2 96376 39816 96376 39816 0 _0636_
rlabel metal3 77112 42952 77112 42952 0 _0637_
rlabel metal2 90888 36344 90888 36344 0 _0638_
rlabel metal2 89488 40376 89488 40376 0 _0639_
rlabel metal3 95872 43848 95872 43848 0 _0640_
rlabel metal3 84448 29512 84448 29512 0 _0641_
rlabel metal3 85848 42616 85848 42616 0 _0642_
rlabel metal3 82600 37240 82600 37240 0 _0643_
rlabel metal2 85848 41832 85848 41832 0 _0644_
rlabel metal2 70336 31864 70336 31864 0 _0645_
rlabel metal3 69160 39032 69160 39032 0 _0646_
rlabel metal3 82824 39592 82824 39592 0 _0647_
rlabel metal3 62328 38136 62328 38136 0 _0648_
rlabel metal2 60032 41160 60032 41160 0 _0649_
rlabel metal2 59976 39256 59976 39256 0 _0650_
rlabel metal3 68824 41160 68824 41160 0 _0651_
rlabel metal2 53032 34496 53032 34496 0 _0652_
rlabel metal3 58184 41160 58184 41160 0 _0653_
rlabel metal2 60200 42672 60200 42672 0 _0654_
rlabel metal2 53368 43344 53368 43344 0 _0655_
rlabel metal2 52248 43568 52248 43568 0 _0656_
rlabel metal3 49168 43512 49168 43512 0 _0657_
rlabel metal3 57120 43624 57120 43624 0 _0658_
rlabel metal2 74760 46312 74760 46312 0 _0659_
rlabel metal3 72296 66136 72296 66136 0 _0660_
rlabel metal2 72296 58660 72296 58660 0 _0661_
rlabel metal2 73080 67032 73080 67032 0 _0662_
rlabel metal2 73752 75992 73752 75992 0 _0663_
rlabel metal2 75432 76048 75432 76048 0 _0664_
rlabel metal2 74648 75824 74648 75824 0 _0665_
rlabel metal3 73024 73976 73024 73976 0 _0666_
rlabel metal2 76048 75096 76048 75096 0 _0667_
rlabel metal3 75656 75656 75656 75656 0 _0668_
rlabel metal2 51240 44716 51240 44716 0 _0669_
rlabel metal2 77560 62776 77560 62776 0 _0670_
rlabel metal3 75936 39592 75936 39592 0 _0671_
rlabel metal3 78232 38024 78232 38024 0 _0672_
rlabel metal3 94528 36680 94528 36680 0 _0673_
rlabel metal2 79016 40040 79016 40040 0 _0674_
rlabel metal3 92568 37352 92568 37352 0 _0675_
rlabel metal2 96432 37464 96432 37464 0 _0676_
rlabel metal2 74648 35280 74648 35280 0 _0677_
rlabel metal2 83944 33600 83944 33600 0 _0678_
rlabel metal2 89432 36288 89432 36288 0 _0679_
rlabel metal3 72352 34328 72352 34328 0 _0680_
rlabel metal3 84952 34888 84952 34888 0 _0681_
rlabel metal2 72408 34888 72408 34888 0 _0682_
rlabel metal3 61096 32760 61096 32760 0 _0683_
rlabel metal2 71904 35112 71904 35112 0 _0684_
rlabel metal3 61712 35672 61712 35672 0 _0685_
rlabel metal3 65408 34216 65408 34216 0 _0686_
rlabel metal3 76888 37352 76888 37352 0 _0687_
rlabel metal2 64624 40600 64624 40600 0 _0688_
rlabel metal3 63840 38808 63840 38808 0 _0689_
rlabel metal3 70504 43512 70504 43512 0 _0690_
rlabel metal3 63000 43736 63000 43736 0 _0691_
rlabel metal2 91672 54320 91672 54320 0 _0692_
rlabel metal3 72464 56280 72464 56280 0 _0693_
rlabel metal2 72520 61824 72520 61824 0 _0694_
rlabel metal2 77280 49000 77280 49000 0 _0695_
rlabel metal2 77672 49616 77672 49616 0 _0696_
rlabel metal3 96600 49896 96600 49896 0 _0697_
rlabel metal2 73640 54096 73640 54096 0 _0698_
rlabel metal2 74592 54264 74592 54264 0 _0699_
rlabel metal2 76216 50288 76216 50288 0 _0700_
rlabel metal2 97496 50008 97496 50008 0 _0701_
rlabel metal3 80640 51464 80640 51464 0 _0702_
rlabel metal3 78904 51464 78904 51464 0 _0703_
rlabel metal2 94808 49784 94808 49784 0 _0704_
rlabel metal2 93296 46872 93296 46872 0 _0705_
rlabel metal2 93296 52024 93296 52024 0 _0706_
rlabel metal2 93240 51072 93240 51072 0 _0707_
rlabel metal3 94864 52136 94864 52136 0 _0708_
rlabel metal2 93688 54320 93688 54320 0 _0709_
rlabel metal2 96376 50176 96376 50176 0 _0710_
rlabel metal2 97384 51912 97384 51912 0 _0711_
rlabel metal2 93408 50792 93408 50792 0 _0712_
rlabel metal2 67928 52136 67928 52136 0 _0713_
rlabel metal2 61040 46536 61040 46536 0 _0714_
rlabel metal2 68712 49112 68712 49112 0 _0715_
rlabel metal2 74312 49168 74312 49168 0 _0716_
rlabel metal3 71120 50008 71120 50008 0 _0717_
rlabel metal2 97496 51520 97496 51520 0 _0718_
rlabel metal2 62216 52304 62216 52304 0 _0719_
rlabel metal3 64232 48328 64232 48328 0 _0720_
rlabel metal3 65576 47208 65576 47208 0 _0721_
rlabel metal3 72800 51352 72800 51352 0 _0722_
rlabel metal2 55160 49392 55160 49392 0 _0723_
rlabel metal3 61376 47992 61376 47992 0 _0724_
rlabel metal2 63448 48216 63448 48216 0 _0725_
rlabel metal2 75152 50344 75152 50344 0 _0726_
rlabel metal2 65128 47208 65128 47208 0 _0727_
rlabel metal2 53144 53032 53144 53032 0 _0728_
rlabel metal2 61768 47936 61768 47936 0 _0729_
rlabel metal3 65240 48216 65240 48216 0 _0730_
rlabel metal2 63952 51128 63952 51128 0 _0731_
rlabel metal2 74648 41104 74648 41104 0 _0732_
rlabel metal2 75320 37520 75320 37520 0 _0733_
rlabel metal2 65688 50120 65688 50120 0 _0734_
rlabel metal3 76384 57736 76384 57736 0 _0735_
rlabel metal2 73752 56952 73752 56952 0 _0736_
rlabel metal3 79688 59192 79688 59192 0 _0737_
rlabel metal2 92792 54712 92792 54712 0 _0738_
rlabel metal2 94752 54712 94752 54712 0 _0739_
rlabel metal2 70168 57456 70168 57456 0 _0740_
rlabel metal2 96488 58184 96488 58184 0 _0741_
rlabel metal2 97608 58800 97608 58800 0 _0742_
rlabel metal2 81592 57288 81592 57288 0 _0743_
rlabel metal3 80136 57736 80136 57736 0 _0744_
rlabel metal2 93072 54712 93072 54712 0 _0745_
rlabel metal3 92568 57736 92568 57736 0 _0746_
rlabel metal3 71456 60760 71456 60760 0 _0747_
rlabel metal3 97720 59864 97720 59864 0 _0748_
rlabel metal3 94752 56616 94752 56616 0 _0749_
rlabel metal3 95032 59304 95032 59304 0 _0750_
rlabel metal2 92232 60256 92232 60256 0 _0751_
rlabel metal3 62272 53704 62272 53704 0 _0752_
rlabel metal2 67424 53704 67424 53704 0 _0753_
rlabel metal3 68656 56056 68656 56056 0 _0754_
rlabel metal2 67592 56280 67592 56280 0 _0755_
rlabel metal2 94584 61096 94584 61096 0 _0756_
rlabel metal2 56728 53872 56728 53872 0 _0757_
rlabel metal2 54488 58464 54488 58464 0 _0758_
rlabel metal2 68040 60256 68040 60256 0 _0759_
rlabel metal3 57120 57064 57120 57064 0 _0760_
rlabel metal3 57512 57736 57512 57736 0 _0761_
rlabel metal2 58968 59696 58968 59696 0 _0762_
rlabel metal2 54376 59024 54376 59024 0 _0763_
rlabel metal2 53144 56616 53144 56616 0 _0764_
rlabel metal2 57400 57456 57400 57456 0 _0765_
rlabel metal3 56448 60200 56448 60200 0 _0766_
rlabel metal2 82040 66864 82040 66864 0 _0767_
rlabel metal3 77672 51352 77672 51352 0 _0768_
rlabel metal2 58520 59416 58520 59416 0 _0769_
rlabel metal3 94528 48888 94528 48888 0 _0770_
rlabel metal3 75152 66248 75152 66248 0 _0771_
rlabel metal2 75768 74424 75768 74424 0 _0772_
rlabel metal2 94024 73640 94024 73640 0 _0773_
rlabel metal2 95928 75208 95928 75208 0 _0774_
rlabel metal3 78960 73528 78960 73528 0 _0775_
rlabel metal3 95088 74760 95088 74760 0 _0776_
rlabel metal2 93408 75096 93408 75096 0 _0777_
rlabel metal3 96432 73304 96432 73304 0 _0778_
rlabel metal2 90888 72968 90888 72968 0 _0779_
rlabel metal2 72296 74704 72296 74704 0 _0780_
rlabel metal3 88872 74872 88872 74872 0 _0781_
rlabel metal2 91448 75152 91448 75152 0 _0782_
rlabel metal2 70056 75768 70056 75768 0 _0783_
rlabel metal3 70168 75096 70168 75096 0 _0784_
rlabel metal3 88984 73304 88984 73304 0 _0785_
rlabel metal3 58800 73976 58800 73976 0 _0786_
rlabel metal3 70672 73864 70672 73864 0 _0787_
rlabel metal3 57232 72744 57232 72744 0 _0788_
rlabel metal3 69048 73976 69048 73976 0 _0789_
rlabel metal2 56448 73976 56448 73976 0 _0790_
rlabel metal3 55832 72408 55832 72408 0 _0791_
rlabel metal2 56280 69496 56280 69496 0 _0792_
rlabel metal2 51408 57848 51408 57848 0 _0793_
rlabel metal3 60368 70056 60368 70056 0 _0794_
rlabel metal2 50232 68880 50232 68880 0 _0795_
rlabel metal2 54600 69328 54600 69328 0 _0796_
rlabel metal2 79464 57960 79464 57960 0 _0797_
rlabel metal2 49784 72240 49784 72240 0 _0798_
rlabel metal2 77280 81704 77280 81704 0 _0799_
rlabel metal2 94584 77336 94584 77336 0 _0800_
rlabel metal3 96992 79576 96992 79576 0 _0801_
rlabel metal2 77896 86352 77896 86352 0 _0802_
rlabel metal2 95256 85176 95256 85176 0 _0803_
rlabel metal3 95704 79688 95704 79688 0 _0804_
rlabel metal2 73920 85736 73920 85736 0 _0805_
rlabel metal2 91224 85904 91224 85904 0 _0806_
rlabel metal2 95200 82152 95200 82152 0 _0807_
rlabel metal2 70616 84392 70616 84392 0 _0808_
rlabel metal2 91224 84392 91224 84392 0 _0809_
rlabel metal2 71960 87192 71960 87192 0 _0810_
rlabel metal2 57904 87640 57904 87640 0 _0811_
rlabel metal3 70000 86520 70000 86520 0 _0812_
rlabel metal2 61600 86632 61600 86632 0 _0813_
rlabel metal2 59752 85512 59752 85512 0 _0814_
rlabel metal2 74760 87024 74760 87024 0 _0815_
rlabel metal2 63784 83048 63784 83048 0 _0816_
rlabel metal2 61544 85624 61544 85624 0 _0817_
rlabel metal2 75320 85512 75320 85512 0 _0818_
rlabel metal2 74872 73416 74872 73416 0 _0819_
rlabel metal2 63504 83720 63504 83720 0 _0820_
rlabel metal2 74984 74312 74984 74312 0 _0821_
rlabel metal2 77560 82768 77560 82768 0 _0822_
rlabel metal2 93240 78876 93240 78876 0 _0823_
rlabel metal3 77504 83384 77504 83384 0 _0824_
rlabel metal2 93352 82824 93352 82824 0 _0825_
rlabel metal3 92848 79352 92848 79352 0 _0826_
rlabel metal2 73192 83384 73192 83384 0 _0827_
rlabel metal3 87360 86856 87360 86856 0 _0828_
rlabel metal2 88312 83888 88312 83888 0 _0829_
rlabel metal2 69720 83776 69720 83776 0 _0830_
rlabel metal2 1848 12432 1848 12432 0 address[0]
rlabel metal3 1302 37464 1302 37464 0 address[1]
rlabel metal3 1302 62440 1302 62440 0 address[2]
rlabel metal3 1246 87416 1246 87416 0 address[3]
rlabel metal3 93184 72408 93184 72408 0 clk
rlabel metal3 86912 72520 86912 72520 0 clknet_0_clk
rlabel metal2 69272 50736 69272 50736 0 clknet_2_0__leaf_clk
rlabel metal2 92008 50176 92008 50176 0 clknet_2_1__leaf_clk
rlabel metal2 52920 76832 52920 76832 0 clknet_2_2__leaf_clk
rlabel metal2 91896 74032 91896 74032 0 clknet_2_3__leaf_clk
rlabel metal2 53816 54992 53816 54992 0 clknet_leaf_0_clk
rlabel metal3 62776 86744 62776 86744 0 clknet_leaf_10_clk
rlabel metal3 62496 74872 62496 74872 0 clknet_leaf_11_clk
rlabel metal2 69496 81984 69496 81984 0 clknet_leaf_12_clk
rlabel metal2 70616 76104 70616 76104 0 clknet_leaf_13_clk
rlabel metal2 67592 75824 67592 75824 0 clknet_leaf_14_clk
rlabel metal2 69608 71400 69608 71400 0 clknet_leaf_15_clk
rlabel metal2 77392 67928 77392 67928 0 clknet_leaf_16_clk
rlabel metal2 81256 74760 81256 74760 0 clknet_leaf_17_clk
rlabel metal3 76776 77224 76776 77224 0 clknet_leaf_18_clk
rlabel metal2 78792 83944 78792 83944 0 clknet_leaf_19_clk
rlabel metal2 64736 53704 64736 53704 0 clknet_leaf_1_clk
rlabel metal2 87696 76664 87696 76664 0 clknet_leaf_20_clk
rlabel metal2 88928 78904 88928 78904 0 clknet_leaf_21_clk
rlabel metal2 90888 88256 90888 88256 0 clknet_leaf_22_clk
rlabel metal3 94136 80360 94136 80360 0 clknet_leaf_23_clk
rlabel metal2 94920 75208 94920 75208 0 clknet_leaf_24_clk
rlabel metal3 92120 74200 92120 74200 0 clknet_leaf_25_clk
rlabel metal3 96208 72520 96208 72520 0 clknet_leaf_26_clk
rlabel metal2 93576 60312 93576 60312 0 clknet_leaf_27_clk
rlabel metal2 91560 66696 91560 66696 0 clknet_leaf_28_clk
rlabel metal2 83496 66976 83496 66976 0 clknet_leaf_29_clk
rlabel metal2 61880 49336 61880 49336 0 clknet_leaf_2_clk
rlabel metal2 86016 54712 86016 54712 0 clknet_leaf_30_clk
rlabel metal2 88200 51016 88200 51016 0 clknet_leaf_31_clk
rlabel metal2 92232 54208 92232 54208 0 clknet_leaf_32_clk
rlabel metal2 98056 53760 98056 53760 0 clknet_leaf_33_clk
rlabel metal2 92008 45416 92008 45416 0 clknet_leaf_34_clk
rlabel metal3 94976 42840 94976 42840 0 clknet_leaf_35_clk
rlabel metal2 94472 34104 94472 34104 0 clknet_leaf_36_clk
rlabel metal2 90888 39928 90888 39928 0 clknet_leaf_38_clk
rlabel metal2 88200 41216 88200 41216 0 clknet_leaf_39_clk
rlabel metal3 62720 55160 62720 55160 0 clknet_leaf_3_clk
rlabel metal2 78792 33712 78792 33712 0 clknet_leaf_40_clk
rlabel metal3 75544 34888 75544 34888 0 clknet_leaf_41_clk
rlabel metal3 77504 45080 77504 45080 0 clknet_leaf_42_clk
rlabel metal3 77728 48216 77728 48216 0 clknet_leaf_43_clk
rlabel metal3 72408 50568 72408 50568 0 clknet_leaf_44_clk
rlabel metal2 66360 43064 66360 43064 0 clknet_leaf_45_clk
rlabel metal2 77224 40040 77224 40040 0 clknet_leaf_46_clk
rlabel metal2 70840 31472 70840 31472 0 clknet_leaf_47_clk
rlabel via2 65352 38024 65352 38024 0 clknet_leaf_48_clk
rlabel metal2 66360 63952 66360 63952 0 clknet_leaf_4_clk
rlabel metal2 54488 33712 54488 33712 0 clknet_leaf_50_clk
rlabel metal3 52808 44072 52808 44072 0 clknet_leaf_51_clk
rlabel metal2 52920 45920 52920 45920 0 clknet_leaf_52_clk
rlabel metal3 64344 70392 64344 70392 0 clknet_leaf_5_clk
rlabel metal3 50120 59976 50120 59976 0 clknet_leaf_6_clk
rlabel metal3 49280 69384 49280 69384 0 clknet_leaf_7_clk
rlabel metal2 49896 76440 49896 76440 0 clknet_leaf_8_clk
rlabel metal2 49560 79968 49560 79968 0 clknet_leaf_9_clk
rlabel metal2 6328 3416 6328 3416 0 data_in[0]
rlabel metal2 18760 3416 18760 3416 0 data_in[1]
rlabel metal2 31192 3416 31192 3416 0 data_in[2]
rlabel metal3 44016 3416 44016 3416 0 data_in[3]
rlabel metal2 56112 3416 56112 3416 0 data_in[4]
rlabel metal2 68824 2856 68824 2856 0 data_in[5]
rlabel metal2 80920 3416 80920 3416 0 data_in[6]
rlabel metal2 93352 3416 93352 3416 0 data_in[7]
rlabel metal2 6776 96376 6776 96376 0 data_out[0]
rlabel metal2 19208 96880 19208 96880 0 data_out[1]
rlabel metal2 31304 97706 31304 97706 0 data_out[2]
rlabel metal2 45080 96376 45080 96376 0 data_out[3]
rlabel metal2 56840 96376 56840 96376 0 data_out[4]
rlabel metal2 68936 96376 68936 96376 0 data_out[5]
rlabel metal2 81368 96880 81368 96880 0 data_out[6]
rlabel metal3 93912 96152 93912 96152 0 data_out[7]
rlabel metal2 73416 52864 73416 52864 0 net1
rlabel metal2 91280 52136 91280 52136 0 net10
rlabel metal2 93688 45640 93688 45640 0 net11
rlabel metal2 75096 45640 75096 45640 0 net12
rlabel metal2 76944 49224 76944 49224 0 net13
rlabel metal3 8120 96040 8120 96040 0 net14
rlabel metal3 24528 95816 24528 95816 0 net15
rlabel metal2 46984 64120 46984 64120 0 net16
rlabel metal2 46312 95816 46312 95816 0 net17
rlabel metal2 57680 96040 57680 96040 0 net18
rlabel metal3 74256 95816 74256 95816 0 net19
rlabel metal2 2184 47488 2184 47488 0 net2
rlabel metal2 88200 73192 88200 73192 0 net20
rlabel metal3 95704 96040 95704 96040 0 net21
rlabel metal2 2184 62832 2184 62832 0 net3
rlabel metal2 68264 61264 68264 61264 0 net4
rlabel metal3 51296 50568 51296 50568 0 net5
rlabel metal2 55384 50624 55384 50624 0 net6
rlabel metal2 31864 3080 31864 3080 0 net7
rlabel metal2 45304 3024 45304 3024 0 net8
rlabel metal2 57064 3136 57064 3136 0 net9
rlabel metal3 50736 55384 50736 55384 0 ram16\[0\].rb.ram1\[0\].rc.mem
rlabel metal3 51744 53480 51744 53480 0 ram16\[0\].rb.ram1\[0\].rc.rd
rlabel metal2 52136 54712 52136 54712 0 ram16\[0\].rb.ram1\[1\].rc.mem
rlabel metal2 52976 54600 52976 54600 0 ram16\[0\].rb.ram1\[1\].rc.rd
rlabel metal2 50008 60760 50008 60760 0 ram16\[0\].rb.ram1\[2\].rc.mem
rlabel metal2 52472 59024 52472 59024 0 ram16\[0\].rb.ram1\[2\].rc.rd
rlabel metal2 67032 67760 67032 67760 0 ram16\[0\].rb.ram1\[3\].rc.mem
rlabel metal1 66472 60200 66472 60200 0 ram16\[0\].rb.ram1\[3\].rc.rd
rlabel metal2 84280 71400 84280 71400 0 ram16\[0\].rb.ram1\[4\].rc.mem
rlabel metal2 85232 50008 85232 50008 0 ram16\[0\].rb.ram1\[4\].rc.rd
rlabel metal2 83888 53928 83888 53928 0 ram16\[0\].rb.ram1\[5\].rc.mem
rlabel metal2 86856 57512 86856 57512 0 ram16\[0\].rb.ram1\[5\].rc.rd
rlabel metal2 84280 45416 84280 45416 0 ram16\[0\].rb.ram1\[6\].rc.mem
rlabel metal2 86296 46256 86296 46256 0 ram16\[0\].rb.ram1\[6\].rc.rd
rlabel metal3 77168 44408 77168 44408 0 ram16\[0\].rb.ram1\[7\].rc.mem
rlabel metal2 80528 44968 80528 44968 0 ram16\[0\].rb.ram1\[7\].rc.rd
rlabel metal3 63896 53144 63896 53144 0 ram16\[10\].rb.ram1\[0\].rc.mem
rlabel metal2 61432 58184 61432 58184 0 ram16\[10\].rb.ram1\[0\].rc.rd
rlabel metal3 64568 56168 64568 56168 0 ram16\[10\].rb.ram1\[1\].rc.mem
rlabel metal3 64120 59080 64120 59080 0 ram16\[10\].rb.ram1\[1\].rc.rd
rlabel metal2 65576 53704 65576 53704 0 ram16\[10\].rb.ram1\[2\].rc.mem
rlabel metal3 65352 58184 65352 58184 0 ram16\[10\].rb.ram1\[2\].rc.rd
rlabel metal2 69496 53144 69496 53144 0 ram16\[10\].rb.ram1\[3\].rc.mem
rlabel metal2 69832 52304 69832 52304 0 ram16\[10\].rb.ram1\[3\].rc.rd
rlabel metal3 92624 56616 92624 56616 0 ram16\[10\].rb.ram1\[4\].rc.mem
rlabel metal2 88704 56728 88704 56728 0 ram16\[10\].rb.ram1\[4\].rc.rd
rlabel metal2 87864 54208 87864 54208 0 ram16\[10\].rb.ram1\[5\].rc.mem
rlabel metal2 86072 52864 86072 52864 0 ram16\[10\].rb.ram1\[5\].rc.rd
rlabel metal2 92232 56616 92232 56616 0 ram16\[10\].rb.ram1\[6\].rc.mem
rlabel metal2 89320 57904 89320 57904 0 ram16\[10\].rb.ram1\[6\].rc.rd
rlabel metal3 79352 53144 79352 53144 0 ram16\[10\].rb.ram1\[7\].rc.mem
rlabel metal2 79016 55216 79016 55216 0 ram16\[10\].rb.ram1\[7\].rc.rd
rlabel metal2 62664 66528 62664 66528 0 ram16\[11\].rb.ram1\[0\].rc.mem
rlabel metal2 61880 61656 61880 61656 0 ram16\[11\].rb.ram1\[0\].rc.rd
rlabel metal3 63616 71064 63616 71064 0 ram16\[11\].rb.ram1\[1\].rc.mem
rlabel metal2 62776 61600 62776 61600 0 ram16\[11\].rb.ram1\[1\].rc.rd
rlabel metal2 63056 73976 63056 73976 0 ram16\[11\].rb.ram1\[2\].rc.mem
rlabel metal3 65968 59864 65968 59864 0 ram16\[11\].rb.ram1\[2\].rc.rd
rlabel metal3 72240 69272 72240 69272 0 ram16\[11\].rb.ram1\[3\].rc.mem
rlabel metal2 70728 52080 70728 52080 0 ram16\[11\].rb.ram1\[3\].rc.rd
rlabel metal2 91000 70448 91000 70448 0 ram16\[11\].rb.ram1\[4\].rc.mem
rlabel metal2 92120 68152 92120 68152 0 ram16\[11\].rb.ram1\[4\].rc.rd
rlabel metal3 95144 69496 95144 69496 0 ram16\[11\].rb.ram1\[5\].rc.mem
rlabel metal3 96152 70056 96152 70056 0 ram16\[11\].rb.ram1\[5\].rc.rd
rlabel metal3 96992 65576 96992 65576 0 ram16\[11\].rb.ram1\[6\].rc.mem
rlabel metal2 93800 65184 93800 65184 0 ram16\[11\].rb.ram1\[6\].rc.rd
rlabel metal3 76160 69272 76160 69272 0 ram16\[11\].rb.ram1\[7\].rc.mem
rlabel metal2 80136 69160 80136 69160 0 ram16\[11\].rb.ram1\[7\].rc.rd
rlabel metal2 51464 37632 51464 37632 0 ram16\[12\].rb.ram1\[0\].rc.mem
rlabel metal2 52192 49112 52192 49112 0 ram16\[12\].rb.ram1\[0\].rc.rd
rlabel metal2 52696 35168 52696 35168 0 ram16\[12\].rb.ram1\[1\].rc.mem
rlabel metal2 53200 50456 53200 50456 0 ram16\[12\].rb.ram1\[1\].rc.rd
rlabel metal2 57400 32984 57400 32984 0 ram16\[12\].rb.ram1\[2\].rc.mem
rlabel metal2 58464 47096 58464 47096 0 ram16\[12\].rb.ram1\[2\].rc.rd
rlabel metal3 68152 32424 68152 32424 0 ram16\[12\].rb.ram1\[3\].rc.mem
rlabel metal2 68264 36008 68264 36008 0 ram16\[12\].rb.ram1\[3\].rc.rd
rlabel metal3 85344 30856 85344 30856 0 ram16\[12\].rb.ram1\[4\].rc.mem
rlabel metal3 87920 47992 87920 47992 0 ram16\[12\].rb.ram1\[4\].rc.rd
rlabel metal2 89544 34160 89544 34160 0 ram16\[12\].rb.ram1\[5\].rc.mem
rlabel metal2 90776 33964 90776 33964 0 ram16\[12\].rb.ram1\[5\].rc.rd
rlabel metal3 96432 34104 96432 34104 0 ram16\[12\].rb.ram1\[6\].rc.mem
rlabel metal2 92736 53032 92736 53032 0 ram16\[12\].rb.ram1\[6\].rc.rd
rlabel metal3 76832 35000 76832 35000 0 ram16\[12\].rb.ram1\[7\].rc.mem
rlabel metal2 77896 33096 77896 33096 0 ram16\[12\].rb.ram1\[7\].rc.rd
rlabel metal2 52472 65464 52472 65464 0 ram16\[13\].rb.ram1\[0\].rc.mem
rlabel metal2 53592 63784 53592 63784 0 ram16\[13\].rb.ram1\[0\].rc.rd
rlabel metal2 51520 64792 51520 64792 0 ram16\[13\].rb.ram1\[1\].rc.mem
rlabel metal2 52472 63840 52472 63840 0 ram16\[13\].rb.ram1\[1\].rc.rd
rlabel metal2 52024 67592 52024 67592 0 ram16\[13\].rb.ram1\[2\].rc.mem
rlabel metal3 57288 66360 57288 66360 0 ram16\[13\].rb.ram1\[2\].rc.rd
rlabel metal3 68768 67704 68768 67704 0 ram16\[13\].rb.ram1\[3\].rc.mem
rlabel metal3 68488 66920 68488 66920 0 ram16\[13\].rb.ram1\[3\].rc.rd
rlabel metal3 88536 69272 88536 69272 0 ram16\[13\].rb.ram1\[4\].rc.mem
rlabel metal2 90216 65744 90216 65744 0 ram16\[13\].rb.ram1\[4\].rc.rd
rlabel metal3 87360 67256 87360 67256 0 ram16\[13\].rb.ram1\[5\].rc.mem
rlabel metal2 90160 66360 90160 66360 0 ram16\[13\].rb.ram1\[5\].rc.rd
rlabel metal2 86072 65688 86072 65688 0 ram16\[13\].rb.ram1\[6\].rc.mem
rlabel metal2 89432 65184 89432 65184 0 ram16\[13\].rb.ram1\[6\].rc.rd
rlabel metal3 79912 66920 79912 66920 0 ram16\[13\].rb.ram1\[7\].rc.mem
rlabel metal2 81480 66192 81480 66192 0 ram16\[13\].rb.ram1\[7\].rc.rd
rlabel metal3 53144 82040 53144 82040 0 ram16\[14\].rb.ram1\[0\].rc.mem
rlabel metal2 59416 78120 59416 78120 0 ram16\[14\].rb.ram1\[0\].rc.rd
rlabel metal2 53592 78820 53592 78820 0 ram16\[14\].rb.ram1\[1\].rc.mem
rlabel metal2 54600 80360 54600 80360 0 ram16\[14\].rb.ram1\[1\].rc.rd
rlabel metal2 53144 80136 53144 80136 0 ram16\[14\].rb.ram1\[2\].rc.mem
rlabel metal2 57064 80360 57064 80360 0 ram16\[14\].rb.ram1\[2\].rc.rd
rlabel metal3 69048 80248 69048 80248 0 ram16\[14\].rb.ram1\[3\].rc.mem
rlabel metal2 70280 79912 70280 79912 0 ram16\[14\].rb.ram1\[3\].rc.rd
rlabel metal2 81368 85904 81368 85904 0 ram16\[14\].rb.ram1\[4\].rc.mem
rlabel metal2 82936 81648 82936 81648 0 ram16\[14\].rb.ram1\[4\].rc.rd
rlabel metal2 82992 83608 82992 83608 0 ram16\[14\].rb.ram1\[5\].rc.mem
rlabel via2 84840 81704 84840 81704 0 ram16\[14\].rb.ram1\[5\].rc.rd
rlabel metal2 81704 80864 81704 80864 0 ram16\[14\].rb.ram1\[6\].rc.mem
rlabel metal3 83720 79464 83720 79464 0 ram16\[14\].rb.ram1\[6\].rc.rd
rlabel metal2 75208 80360 75208 80360 0 ram16\[14\].rb.ram1\[7\].rc.mem
rlabel metal2 76216 78344 76216 78344 0 ram16\[14\].rb.ram1\[7\].rc.rd
rlabel metal2 55160 75264 55160 75264 0 ram16\[15\].rb.ram1\[0\].rc.mem
rlabel metal3 59080 78008 59080 78008 0 ram16\[15\].rb.ram1\[0\].rc.rd
rlabel metal2 53592 75656 53592 75656 0 ram16\[15\].rb.ram1\[1\].rc.mem
rlabel metal2 57288 77392 57288 77392 0 ram16\[15\].rb.ram1\[1\].rc.rd
rlabel metal2 52920 74872 52920 74872 0 ram16\[15\].rb.ram1\[2\].rc.mem
rlabel metal2 56616 76944 56616 76944 0 ram16\[15\].rb.ram1\[2\].rc.rd
rlabel metal2 66696 76160 66696 76160 0 ram16\[15\].rb.ram1\[3\].rc.mem
rlabel metal2 67256 79240 67256 79240 0 ram16\[15\].rb.ram1\[3\].rc.rd
rlabel metal2 81928 76160 81928 76160 0 ram16\[15\].rb.ram1\[4\].rc.mem
rlabel metal3 84392 78792 84392 78792 0 ram16\[15\].rb.ram1\[4\].rc.rd
rlabel metal2 85400 75936 85400 75936 0 ram16\[15\].rb.ram1\[5\].rc.mem
rlabel metal3 85232 79576 85232 79576 0 ram16\[15\].rb.ram1\[5\].rc.rd
rlabel metal2 84616 74760 84616 74760 0 ram16\[15\].rb.ram1\[6\].rc.mem
rlabel metal2 85288 77280 85288 77280 0 ram16\[15\].rb.ram1\[6\].rc.rd
rlabel metal2 76104 75936 76104 75936 0 ram16\[15\].rb.ram1\[7\].rc.mem
rlabel metal3 77448 78008 77448 78008 0 ram16\[15\].rb.ram1\[7\].rc.rd
rlabel metal2 51912 44044 51912 44044 0 ram16\[1\].rb.ram1\[0\].rc.mem
rlabel metal2 52976 44968 52976 44968 0 ram16\[1\].rb.ram1\[0\].rc.rd
rlabel metal3 59192 42840 59192 42840 0 ram16\[1\].rb.ram1\[1\].rc.mem
rlabel metal2 59752 50736 59752 50736 0 ram16\[1\].rb.ram1\[1\].rc.rd
rlabel metal2 62552 39088 62552 39088 0 ram16\[1\].rb.ram1\[2\].rc.mem
rlabel metal2 62552 51240 62552 51240 0 ram16\[1\].rb.ram1\[2\].rc.rd
rlabel metal2 70280 40992 70280 40992 0 ram16\[1\].rb.ram1\[3\].rc.mem
rlabel metal2 70448 50568 70448 50568 0 ram16\[1\].rb.ram1\[3\].rc.rd
rlabel metal3 83944 38136 83944 38136 0 ram16\[1\].rb.ram1\[4\].rc.mem
rlabel metal2 85400 49672 85400 49672 0 ram16\[1\].rb.ram1\[4\].rc.rd
rlabel metal3 87976 42728 87976 42728 0 ram16\[1\].rb.ram1\[5\].rc.mem
rlabel metal2 87528 50120 87528 50120 0 ram16\[1\].rb.ram1\[5\].rc.rd
rlabel metal2 96040 40264 96040 40264 0 ram16\[1\].rb.ram1\[6\].rc.mem
rlabel metal2 94920 44912 94920 44912 0 ram16\[1\].rb.ram1\[6\].rc.rd
rlabel metal2 77784 43344 77784 43344 0 ram16\[1\].rb.ram1\[7\].rc.mem
rlabel metal2 79800 43400 79800 43400 0 ram16\[1\].rb.ram1\[7\].rc.rd
rlabel metal2 64232 41104 64232 41104 0 ram16\[2\].rb.ram1\[0\].rc.mem
rlabel metal2 65912 60592 65912 60592 0 ram16\[2\].rb.ram1\[0\].rc.rd
rlabel metal2 62776 35840 62776 35840 0 ram16\[2\].rb.ram1\[1\].rc.mem
rlabel metal2 64344 37800 64344 37800 0 ram16\[2\].rb.ram1\[1\].rc.rd
rlabel metal3 62944 33992 62944 33992 0 ram16\[2\].rb.ram1\[2\].rc.mem
rlabel metal3 63952 34328 63952 34328 0 ram16\[2\].rb.ram1\[2\].rc.rd
rlabel metal2 72632 34160 72632 34160 0 ram16\[2\].rb.ram1\[3\].rc.mem
rlabel metal2 72744 52136 72744 52136 0 ram16\[2\].rb.ram1\[3\].rc.rd
rlabel metal2 85960 34944 85960 34944 0 ram16\[2\].rb.ram1\[4\].rc.mem
rlabel metal3 87920 36568 87920 36568 0 ram16\[2\].rb.ram1\[4\].rc.rd
rlabel metal2 89544 37296 89544 37296 0 ram16\[2\].rb.ram1\[5\].rc.mem
rlabel metal2 90440 51184 90440 51184 0 ram16\[2\].rb.ram1\[5\].rc.rd
rlabel metal3 96824 37240 96824 37240 0 ram16\[2\].rb.ram1\[6\].rc.mem
rlabel metal3 96600 39704 96600 39704 0 ram16\[2\].rb.ram1\[6\].rc.rd
rlabel metal3 77000 38696 77000 38696 0 ram16\[2\].rb.ram1\[7\].rc.mem
rlabel metal3 82152 39704 82152 39704 0 ram16\[2\].rb.ram1\[7\].rc.rd
rlabel metal2 64288 45976 64288 45976 0 ram16\[3\].rb.ram1\[0\].rc.mem
rlabel metal2 66024 50736 66024 50736 0 ram16\[3\].rb.ram1\[0\].rc.rd
rlabel metal2 64344 46648 64344 46648 0 ram16\[3\].rb.ram1\[1\].rc.mem
rlabel metal2 64064 51576 64064 51576 0 ram16\[3\].rb.ram1\[1\].rc.rd
rlabel metal2 66472 46088 66472 46088 0 ram16\[3\].rb.ram1\[2\].rc.mem
rlabel metal2 63616 59976 63616 59976 0 ram16\[3\].rb.ram1\[2\].rc.rd
rlabel metal2 71624 48216 71624 48216 0 ram16\[3\].rb.ram1\[3\].rc.mem
rlabel metal3 72800 51464 72800 51464 0 ram16\[3\].rb.ram1\[3\].rc.rd
rlabel metal2 97832 51296 97832 51296 0 ram16\[3\].rb.ram1\[4\].rc.mem
rlabel metal2 94864 52248 94864 52248 0 ram16\[3\].rb.ram1\[4\].rc.rd
rlabel metal2 96488 48216 96488 48216 0 ram16\[3\].rb.ram1\[5\].rc.mem
rlabel via2 91224 50008 91224 50008 0 ram16\[3\].rb.ram1\[5\].rc.rd
rlabel metal2 96264 47544 96264 47544 0 ram16\[3\].rb.ram1\[6\].rc.mem
rlabel metal2 92624 52808 92624 52808 0 ram16\[3\].rb.ram1\[6\].rc.rd
rlabel metal3 79856 49672 79856 49672 0 ram16\[3\].rb.ram1\[7\].rc.mem
rlabel metal3 83048 59976 83048 59976 0 ram16\[3\].rb.ram1\[7\].rc.rd
rlabel metal3 56952 56728 56952 56728 0 ram16\[4\].rb.ram1\[0\].rc.mem
rlabel metal2 56616 60536 56616 60536 0 ram16\[4\].rb.ram1\[0\].rc.rd
rlabel metal3 57400 56616 57400 56616 0 ram16\[4\].rb.ram1\[1\].rc.mem
rlabel metal3 57064 59864 57064 59864 0 ram16\[4\].rb.ram1\[1\].rc.rd
rlabel metal2 56784 57512 56784 57512 0 ram16\[4\].rb.ram1\[2\].rc.mem
rlabel metal3 59472 59864 59472 59864 0 ram16\[4\].rb.ram1\[2\].rc.rd
rlabel metal2 68544 54376 68544 54376 0 ram16\[4\].rb.ram1\[3\].rc.mem
rlabel metal2 69328 60984 69328 60984 0 ram16\[4\].rb.ram1\[3\].rc.rd
rlabel metal2 96488 57568 96488 57568 0 ram16\[4\].rb.ram1\[4\].rc.mem
rlabel metal2 95032 63056 95032 63056 0 ram16\[4\].rb.ram1\[4\].rc.rd
rlabel metal2 97160 57344 97160 57344 0 ram16\[4\].rb.ram1\[5\].rc.mem
rlabel metal3 95648 62888 95648 62888 0 ram16\[4\].rb.ram1\[5\].rc.rd
rlabel metal2 96880 56616 96880 56616 0 ram16\[4\].rb.ram1\[6\].rc.mem
rlabel metal2 96432 60088 96432 60088 0 ram16\[4\].rb.ram1\[6\].rc.rd
rlabel metal3 80864 56952 80864 56952 0 ram16\[4\].rb.ram1\[7\].rc.mem
rlabel metal2 82376 62636 82376 62636 0 ram16\[4\].rb.ram1\[7\].rc.rd
rlabel metal2 51688 69888 51688 69888 0 ram16\[5\].rb.ram1\[0\].rc.mem
rlabel metal2 52920 63672 52920 63672 0 ram16\[5\].rb.ram1\[0\].rc.rd
rlabel metal3 57624 71624 57624 71624 0 ram16\[5\].rb.ram1\[1\].rc.mem
rlabel metal3 56112 69496 56112 69496 0 ram16\[5\].rb.ram1\[1\].rc.rd
rlabel metal3 58744 71064 58744 71064 0 ram16\[5\].rb.ram1\[2\].rc.mem
rlabel metal2 59976 69608 59976 69608 0 ram16\[5\].rb.ram1\[2\].rc.rd
rlabel metal2 71512 74480 71512 74480 0 ram16\[5\].rb.ram1\[3\].rc.mem
rlabel metal2 69888 74760 69888 74760 0 ram16\[5\].rb.ram1\[3\].rc.rd
rlabel metal2 90552 73808 90552 73808 0 ram16\[5\].rb.ram1\[4\].rc.mem
rlabel metal2 90552 71008 90552 71008 0 ram16\[5\].rb.ram1\[4\].rc.rd
rlabel metal3 93352 74984 93352 74984 0 ram16\[5\].rb.ram1\[5\].rc.mem
rlabel metal2 91672 74648 91672 74648 0 ram16\[5\].rb.ram1\[5\].rc.rd
rlabel metal3 97104 74200 97104 74200 0 ram16\[5\].rb.ram1\[6\].rc.mem
rlabel metal2 94920 71400 94920 71400 0 ram16\[5\].rb.ram1\[6\].rc.rd
rlabel metal3 76608 73192 76608 73192 0 ram16\[5\].rb.ram1\[7\].rc.mem
rlabel metal2 81592 63168 81592 63168 0 ram16\[5\].rb.ram1\[7\].rc.rd
rlabel metal2 67256 85400 67256 85400 0 ram16\[6\].rb.ram1\[0\].rc.mem
rlabel metal2 62272 78008 62272 78008 0 ram16\[6\].rb.ram1\[0\].rc.rd
rlabel metal2 62776 87416 62776 87416 0 ram16\[6\].rb.ram1\[1\].rc.mem
rlabel metal3 61376 78792 61376 78792 0 ram16\[6\].rb.ram1\[1\].rc.rd
rlabel metal2 59304 86520 59304 86520 0 ram16\[6\].rb.ram1\[2\].rc.mem
rlabel metal2 60424 85512 60424 85512 0 ram16\[6\].rb.ram1\[2\].rc.rd
rlabel metal2 72296 87024 72296 87024 0 ram16\[6\].rb.ram1\[3\].rc.mem
rlabel metal2 70616 80976 70616 80976 0 ram16\[6\].rb.ram1\[3\].rc.rd
rlabel metal3 93072 84952 93072 84952 0 ram16\[6\].rb.ram1\[4\].rc.mem
rlabel metal2 90776 83832 90776 83832 0 ram16\[6\].rb.ram1\[4\].rc.rd
rlabel metal3 97104 84392 97104 84392 0 ram16\[6\].rb.ram1\[5\].rc.mem
rlabel metal2 95592 81872 95592 81872 0 ram16\[6\].rb.ram1\[5\].rc.rd
rlabel metal2 96152 80920 96152 80920 0 ram16\[6\].rb.ram1\[6\].rc.mem
rlabel metal2 97832 78736 97832 78736 0 ram16\[6\].rb.ram1\[6\].rc.rd
rlabel metal3 76776 85736 76776 85736 0 ram16\[6\].rb.ram1\[7\].rc.mem
rlabel metal2 80304 78008 80304 78008 0 ram16\[6\].rb.ram1\[7\].rc.rd
rlabel metal2 62888 79688 62888 79688 0 ram16\[7\].rb.ram1\[0\].rc.mem
rlabel metal2 63448 80808 63448 80808 0 ram16\[7\].rb.ram1\[0\].rc.rd
rlabel metal3 58408 85176 58408 85176 0 ram16\[7\].rb.ram1\[1\].rc.mem
rlabel metal2 59192 78792 59192 78792 0 ram16\[7\].rb.ram1\[1\].rc.rd
rlabel metal2 54432 86520 54432 86520 0 ram16\[7\].rb.ram1\[2\].rc.mem
rlabel metal2 54040 85848 54040 85848 0 ram16\[7\].rb.ram1\[2\].rc.rd
rlabel metal2 70392 86464 70392 86464 0 ram16\[7\].rb.ram1\[3\].rc.mem
rlabel metal2 69272 83216 69272 83216 0 ram16\[7\].rb.ram1\[3\].rc.rd
rlabel metal3 89264 86520 89264 86520 0 ram16\[7\].rb.ram1\[4\].rc.mem
rlabel metal3 87864 85176 87864 85176 0 ram16\[7\].rb.ram1\[4\].rc.rd
rlabel metal3 92904 84168 92904 84168 0 ram16\[7\].rb.ram1\[5\].rc.mem
rlabel metal3 87136 83720 87136 83720 0 ram16\[7\].rb.ram1\[5\].rc.rd
rlabel metal3 93184 79688 93184 79688 0 ram16\[7\].rb.ram1\[6\].rc.mem
rlabel metal2 94360 79128 94360 79128 0 ram16\[7\].rb.ram1\[6\].rc.rd
rlabel metal2 76440 84112 76440 84112 0 ram16\[7\].rb.ram1\[7\].rc.mem
rlabel metal2 78344 81648 78344 81648 0 ram16\[7\].rb.ram1\[7\].rc.rd
rlabel metal3 52976 41832 52976 41832 0 ram16\[8\].rb.ram1\[0\].rc.mem
rlabel metal2 54600 51352 54600 51352 0 ram16\[8\].rb.ram1\[0\].rc.rd
rlabel metal2 56728 39088 56728 39088 0 ram16\[8\].rb.ram1\[1\].rc.mem
rlabel metal3 57624 50680 57624 50680 0 ram16\[8\].rb.ram1\[1\].rc.rd
rlabel metal3 58128 35448 58128 35448 0 ram16\[8\].rb.ram1\[2\].rc.mem
rlabel metal3 62104 51240 62104 51240 0 ram16\[8\].rb.ram1\[2\].rc.rd
rlabel metal2 69608 37576 69608 37576 0 ram16\[8\].rb.ram1\[3\].rc.mem
rlabel metal2 69776 50568 69776 50568 0 ram16\[8\].rb.ram1\[3\].rc.rd
rlabel metal2 82152 34216 82152 34216 0 ram16\[8\].rb.ram1\[4\].rc.mem
rlabel metal2 81368 49224 81368 49224 0 ram16\[8\].rb.ram1\[4\].rc.rd
rlabel metal2 90664 41216 90664 41216 0 ram16\[8\].rb.ram1\[5\].rc.mem
rlabel metal2 84448 48552 84448 48552 0 ram16\[8\].rb.ram1\[5\].rc.rd
rlabel metal3 92792 44296 92792 44296 0 ram16\[8\].rb.ram1\[6\].rc.mem
rlabel metal2 91224 45024 91224 45024 0 ram16\[8\].rb.ram1\[6\].rc.rd
rlabel metal2 75208 38976 75208 38976 0 ram16\[8\].rb.ram1\[7\].rc.mem
rlabel metal2 77336 47880 77336 47880 0 ram16\[8\].rb.ram1\[7\].rc.rd
rlabel metal2 52248 47936 52248 47936 0 ram16\[9\].rb.ram1\[0\].rc.mem
rlabel metal2 54376 48944 54376 48944 0 ram16\[9\].rb.ram1\[0\].rc.rd
rlabel metal2 53592 47488 53592 47488 0 ram16\[9\].rb.ram1\[1\].rc.mem
rlabel metal2 54376 50456 54376 50456 0 ram16\[9\].rb.ram1\[1\].rc.rd
rlabel metal2 58296 46536 58296 46536 0 ram16\[9\].rb.ram1\[2\].rc.mem
rlabel metal2 58744 50232 58744 50232 0 ram16\[9\].rb.ram1\[2\].rc.rd
rlabel metal2 69832 45472 69832 45472 0 ram16\[9\].rb.ram1\[3\].rc.mem
rlabel metal3 69216 58520 69216 58520 0 ram16\[9\].rb.ram1\[3\].rc.rd
rlabel metal2 92232 48216 92232 48216 0 ram16\[9\].rb.ram1\[4\].rc.mem
rlabel metal2 83832 49336 83832 49336 0 ram16\[9\].rb.ram1\[4\].rc.rd
rlabel metal3 91560 47544 91560 47544 0 ram16\[9\].rb.ram1\[5\].rc.mem
rlabel metal2 86296 49672 86296 49672 0 ram16\[9\].rb.ram1\[5\].rc.rd
rlabel metal3 91672 45752 91672 45752 0 ram16\[9\].rb.ram1\[6\].rc.mem
rlabel metal3 86632 47432 86632 47432 0 ram16\[9\].rb.ram1\[6\].rc.rd
rlabel metal2 75656 47208 75656 47208 0 ram16\[9\].rb.ram1\[7\].rc.mem
rlabel metal2 78120 48160 78120 48160 0 ram16\[9\].rb.ram1\[7\].rc.rd
rlabel metal3 95816 25144 95816 25144 0 rd_wr
<< properties >>
string FIXED_BBOX 0 0 100000 100000
<< end >>
